netcdf ukcp18-land-prob-uk-25km-all {
dimensions:
	time = UNLIMITED ; // (12 currently)
	bnds = 2 ;
	projection_y_coordinate = 52 ;
	projection_x_coordinate = 39 ;
variables:
	double climatology_bounds(time, bnds) ;
	float example_var(time, projection_y_coordinate, projection_x_coordinate) ;
		example_var:_FillValue = 1.e+20f ;
		example_var:standard_name = "air_temperature" ;
		example_var:long_name = "Monthly mean air temperature" ;
		example_var:units = "degC" ;
		example_var:cell_methods = "time: mid_range within days time: mean over days" ;
		example_var:coordinates = "latitude longitude" ;
		example_var:grid_mapping = "transverse_mercator" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	double time_bnds(time, bnds) ;
	double latitude(projection_y_coordinate, projection_x_coordinate) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:grid_mapping = "transverse_mercator" ;
	double longitude(projection_y_coordinate, projection_x_coordinate) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
		longitude:grid_mapping = "transverse_mercator" ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	double time(time) ;
		time:axis = "T" ;
		time:units = "hours since 1851-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "standard" ;
		time:climatology = "climatology_bounds" ;
	int season_year(time) ;
		season_year:units = "1" ;
		season_year:long_name = "season_year" ;

// global attributes:
		:comment = "These data are part of the test suite for the data-factory." ;
		:references = "" ;
		:short_name = "temp data" ;
		:source = "a project" ;
		:title = "Great data at your service" ;
		:Conventions = "CF-1.5" ;
		:history = "Wed Sep 13 08:47:03 2017: ncks -d projection_x_coordinate,,,5 -d projection_y_coordinate,,,5 -v example_var osgb_5km.nc osgb_25km.nc" ;
		:NCO = "\"4.5.5\"" ;
data:

 climatology_bounds =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 example_var =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.815, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 273.7442, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.5787, 276.6121, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.923, 276.0981, 274.9792, 
    274.7773, 275.5051, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.5666, 275.8101, 
    275.2739, 275.3267, 274.6761, 273.4642, 273.7743, 273.6353, 276.8704, 
    274.9566, 272.5102, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.197, 275.3978, 
    275.0655, 275.0132, 274.683, 274.3341, 274.0203, 273.8073, 274.0299, 
    273.7935, 273.3065, 272.8606, 272.8433, 272.9532, 273.8348, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.8535, 275.7036, 
    275.2146, 274.5898, 274.358, 274.3236, 274.12, 274.0012, 273.8219, 
    273.8803, 273.6188, 273.4129, 273.258, 273.1212, 273.6964, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 272.6061, 
    274.3033, 274.2682, 274.1063, 273.7565, 273.594, 273.4839, 273.5007, 
    273.3772, 273.4059, 273.4758, 273.6457, 274.1679, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.6629, 273.664, 
    273.8607, 274.1182, 274.1404, 273.9467, 273.7168, 273.5708, 273.41, 
    273.3702, 273.4179, 273.4111, 273.4821, 273.7307, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.3188, 275.8051, 274.6164, 
    274.2485, 273.8336, 274.1509, 274.1849, 274.0236, 273.7517, 273.4882, 
    273.4241, 273.3399, 273.265, 273.2482, 273.3008, 273.3338, 273.5894, 
    274.674, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.3584, 276.6918, 275.5082, 
    274.4218, 273.6973, 273.7725, 273.8806, 273.7125, 273.6548, 273.3058, 
    273.2671, 273.183, 273.1735, 273.1343, 273.206, 273.1852, 273.2312, 
    273.6894, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.6248, 273.6552, 
    273.61, 273.763, 273.6457, 273.5505, 273.2955, 273.1315, 273.0113, 
    273.0928, 273.1564, 273.1323, 273.0802, 273.1141, 273.5402, 274.1198, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.066, 273.5825, 
    273.5178, 273.5542, 273.5267, 273.406, 273.2063, 273.0175, 272.9144, 
    273.0118, 273.1045, 273.0795, 273.0966, 273.2356, 273.5695, 274.0573, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.9515, 273.3854, 
    273.6091, 273.7908, 273.495, 273.1366, 273.0495, 272.9431, 272.9258, 
    273.0065, 273.0722, 273.2086, 273.4518, 273.6045, 273.8661, 274.4095, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.9178, 274.0201, 
    273.2295, 273.6597, 273.5202, 273.2575, 272.6971, 272.8023, 272.7757, 
    272.9611, 273.0713, 273.1576, 273.5469, 273.8129, 274.164, 274.6833, 
    273.6326, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.3962, 273.7864, 
    273.6519, 273.4306, 273.0176, 272.5983, 272.6927, 272.8017, 272.993, 
    273.0954, 273.213, 273.7189, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.3289, _, _, 
    274.2908, 273.4806, 272.8439, 272.619, 272.6922, 272.9311, 273.0877, 
    273.1241, 273.3505, 273.7775, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 272.9259, 
    272.8, 272.5684, 272.7168, 273.0655, 273.1351, 273.1459, 273.5427, 
    274.2561, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.2362, 
    272.6408, 272.4566, 272.5643, 273.1471, 273.1637, 273.1833, 273.7289, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.7384, 
    272.4114, 272.2245, 272.5965, 273.094, 273.1198, 273.3903, 273.842, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 275.6613, 275.4386, 275.3081, 274.8506, 
    274.6239, 275.6245, _, _, 275.3608, _, _, 271.2096, 271.9632, 272.1688, 
    272.1529, 272.7043, 272.9209, 273.0388, 273.709, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 275.6014, 275.5528, 275.2434, 275.3192, 275.1284, 
    274.9224, 275.673, _, _, _, _, _, 272.9792, 272.4477, 271.8863, 272.1363, 
    272.7928, 273.2805, 273.6632, 274.2382, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 275.4948, 275.334, 275.1112, 275.2243, 275.2239, 
    275.1408, 275.5385, _, _, _, _, _, 272.364, 272.3522, 272.0014, 272.382, 
    272.9294, 273.6098, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 275.625, 275.4246, 275.446, 275.3289, 275.5323, 
    272.929, _, 272.6642, 272.8083, 273.0244, 272.6112, 272.416, 272.3616, 
    272.3127, 272.6352, 273.2651, 273.6307, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, 276.0988, 276.2626, 275.5751, 276.1894, _, _, 
    273.7885, 272.9677, 272.9892, 272.9733, 272.7492, 272.5034, 272.4246, 
    272.6842, 273.3778, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 272.4972, _, _, 273.0905, 
    272.5799, 272.2873, 272.2141, 272.4607, 272.5124, 272.8705, 273.681, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.6299, 273.8045, 272.9554, 
    273.016, 272.582, 272.5377, 272.5464, 272.5364, 272.7685, 273.4315, 
    274.1588, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 275.9141, _, 273.7515, 273.2482, 
    272.8162, 272.5772, 272.5859, 272.7245, 272.982, 273.4571, 273.7173, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 272.64, 272.6273, 272.5819, 
    272.3626, 272.5283, 272.8858, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.1064, 273.2414, 272.8363, 
    271.8817, 271.7217, 272.0031, 272.3787, 272.5001, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 275.7136, 272.8887, 273.6316, 
    272.4091, 271.5261, 271.3341, 271.5186, 271.8918, 272.1831, 273.798, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 272.3977, 273.6611, 272.2593, 
    271.4695, 271.2054, 271.1317, 271.513, 271.7739, 272.1605, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 272.8413, 271.874, 272.0689, 
    271.7602, 271.2846, 270.9272, 271.5122, 272.2455, 272.968, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.1317, 273.3142, 272.3943, 
    272.1693, 272.1148, 272.1014, 272.1369, 272.2214, 272.5063, 273.0525, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 273.4163, _, 273.7289, 274.7257, 273.8685, 
    272.8776, 272.4667, 272.5556, 272.7847, 273.111, 273.2295, 273.2376, 
    273.4833, 277.2598, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 274.75, _, 275.5195, _, 273.9503, 
    273.6555, 272.5886, 272.5676, 273.0975, 273.7679, 275.7294, 274.2314, 
    274.0469, 272.6303, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 274.633, 275.6437, _, _, 275.0587, 
    274.4641, 272.9795, 272.5568, 274.3294, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 272.9502, 272.671, _, _, 275.5395, 
    273.8679, 272.8385, 272.6452, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 272.7166, 275.6907, _, _, 275.8782, 
    273.9153, 273.5312, 273.3106, 273.2072, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.742, 273.6766, 
    274.1006, 274.295, 273.9938, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.5934, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.4048, 
    274.6864, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    275.4346, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    273.8993, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    273.7964, 273.4259, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.4728, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 274.427, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.3273, 276.6361, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.7787, 276.0304, 275.3383, 
    275.5166, 276.214, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.2371, 275.5266, 
    275.0324, 275.3406, 276.0994, 274.2108, 274.1145, 274.2551, 276.3387, 
    274.9136, 273.2253, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.8929, 275.1852, 
    274.9364, 275.0041, 274.762, 274.544, 274.3734, 274.4084, 274.7926, 
    274.7022, 274.4137, 274.004, 274.0634, 274.3484, 274.5789, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.7339, 275.6283, 
    275.2116, 274.7502, 274.6407, 274.4118, 274.385, 274.6836, 274.8198, 
    274.9934, 274.7333, 274.6384, 274.6424, 274.7417, 275.2556, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.1646, 
    274.4049, 274.5711, 274.2708, 273.9138, 274.1301, 274.4152, 274.7047, 
    274.5583, 274.6941, 274.9213, 275.2301, 275.6255, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.5486, 273.7276, 
    273.7892, 274.2621, 274.4492, 274.1509, 273.8976, 274.1331, 274.3804, 
    274.6083, 274.7102, 274.7742, 275.0374, 275.4354, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.9236, 275.7664, 274.9266, 
    274.4267, 273.9111, 274.2296, 274.4073, 274.3988, 274.0713, 273.8517, 
    274.1232, 274.4696, 274.6086, 274.5849, 274.7056, 274.9595, 275.3991, 
    275.0602, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.5524, 276.1527, 275.3986, 
    274.5336, 273.7316, 273.8499, 274.1237, 274.2268, 274.3573, 274.004, 
    274.2351, 274.4793, 274.6279, 274.5158, 274.67, 274.8852, 275.0754, 
    275.4918, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.7601, 273.8406, 
    273.8639, 274.1677, 274.3431, 274.6237, 274.444, 274.3478, 274.3908, 
    274.6204, 274.7084, 274.7513, 274.886, 274.9793, 275.3075, 275.8022, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.3671, 273.943, 
    273.9407, 274.1035, 274.4405, 274.6407, 274.5475, 274.3716, 274.3226, 
    274.5454, 274.7052, 274.7894, 274.9027, 275.0377, 275.3265, 275.7375, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.3681, 273.8561, 
    274.1381, 274.5875, 274.6662, 274.4664, 274.3563, 274.1379, 274.3036, 
    274.5181, 274.6822, 274.9113, 275.1432, 275.2476, 275.4861, 275.9287, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.5699, 274.4461, 
    273.6741, 274.2279, 274.5779, 274.6217, 274.0834, 274.043, 273.9734, 
    274.3375, 274.5504, 274.7538, 275.2389, 275.4324, 275.7144, 276.0663, 
    275.3051, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.7876, 274.2406, 
    274.3954, 274.6064, 274.4594, 273.9572, 273.9295, 274.0694, 274.3463, 
    274.544, 274.8076, 275.3871, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.587, _, _, 275.1716, 
    274.8085, 274.3193, 273.9691, 273.921, 274.1462, 274.3811, 274.5319, 
    274.9171, 275.4264, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.4341, 
    274.2449, 273.8823, 273.9, 274.2332, 274.4022, 274.555, 275.1704, 
    275.8835, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.4829, 
    274.1206, 273.7549, 273.7157, 274.291, 274.4492, 274.584, 275.3736, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.5911, 
    273.8515, 273.6032, 273.8953, 274.3239, 274.4208, 274.7993, 275.4044, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 275.3522, 275.3269, 275.3515, 275.1971, 
    275.1561, 276.1053, _, _, 276.1626, _, _, 273.3275, 273.5982, 273.6083, 
    273.5418, 274.0356, 274.2252, 274.263, 275.0761, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 275.3501, 275.3593, 275.2289, 275.4401, 275.4267, 
    275.3355, 276.1306, _, _, _, _, _, 274.1703, 273.9329, 273.3785, 
    273.3687, 274.1692, 274.7525, 274.95, 275.6091, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 275.3582, 275.2535, 275.1436, 275.3851, 275.5177, 
    275.5742, 276.0385, _, _, _, _, _, 273.9767, 273.9096, 273.4521, 
    273.4686, 274.388, 275.2178, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 275.5432, 275.464, 275.6378, 275.6408, 275.9878, 
    274.5434, _, 273.4655, 273.7004, 273.7882, 273.6934, 273.8969, 273.9327, 
    273.7212, 273.9047, 274.8221, 275.3414, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, 276.0825, 276.4227, 275.8899, 276.5591, _, _, 
    274.1661, 273.8936, 273.8502, 273.8794, 273.9103, 273.9805, 273.7927, 
    274.076, 275.0172, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.4655, _, _, 273.9453, 
    273.6717, 273.5397, 273.5766, 273.8699, 273.9074, 274.2567, 275.2686, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.0529, 274.6146, 274.1128, 
    273.8799, 273.7227, 273.7419, 273.8132, 273.8943, 274.1922, 274.904, 
    275.6499, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 276.0593, _, 274.5692, 274.0592, 
    273.759, 273.7346, 273.8499, 274.0665, 274.3382, 274.8474, 275.7321, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.7586, 273.606, 273.5797, 
    273.4709, 273.8598, 274.3505, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.4992, 274.0927, 273.7041, 
    272.8015, 272.678, 273.0527, 273.5929, 274.0648, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 276.2303, 274.6797, 274.2361, 
    273.2683, 272.2988, 272.2135, 272.5798, 273.0887, 273.5007, 274.8781, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 273.9469, 274.0688, 272.817, 
    272.0021, 271.8547, 271.998, 272.686, 273.2383, 273.5464, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 274.4148, 272.327, 272.2107, 
    272.4168, 271.9186, 271.5723, 272.1366, 273.2629, 274.3461, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.6241, 274.0187, 272.8925, 
    272.6013, 272.6739, 272.6631, 272.6409, 272.7848, 273.3787, 274.459, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 273.6962, _, 275.3633, 274.8044, 274.3253, 
    273.3923, 272.9263, 272.9264, 273.1856, 273.6246, 273.8449, 274.1813, 
    274.8162, 277.2619, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 274.791, _, 275.649, _, 275.5231, 
    273.9615, 273.2611, 273.2097, 273.7442, 274.5295, 275.6678, 275.2564, 
    275.3631, 274.3575, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 275.9871, 275.6747, _, _, 275.8714, 
    274.4156, 273.6244, 273.484, 275.9219, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 274.1632, 274.0499, _, _, 275.4635, 
    274.3759, 273.8443, 274.1181, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 274.6932, 275.7061, _, _, 276.0888, 
    274.4311, 274.3372, 274.5145, 274.7378, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.8929, 275.3738, 
    275.1476, 275.6245, 274.1898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.0532, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.691, 
    276.0789, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.6397, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    275.2664, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    275.4496, 275.5771, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.8039, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 278.1825, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.0133, 280.735, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.3424, 280.6591, 280.2848, 
    279.741, 280.4755, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.4836, 279.9595, 
    279.7771, 280.3055, 280.134, 280.1389, 280.2509, 280.1672, 280.5324, 
    280.2654, 280.327, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.3196, 279.9873, 
    279.9673, 280.2491, 280.3081, 280.2103, 280.1155, 280.1479, 280.0893, 
    280.0542, 280.0735, 279.9821, 279.944, 279.9792, 275.9931, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.3687, 280.3643, 
    280.3302, 280.3434, 280.1249, 280.0952, 280.1382, 280.142, 279.9579, 
    280.0583, 279.9921, 280.006, 280.0464, 280.0282, 280.0791, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.3313, 
    280.4711, 280.1763, 280.1446, 279.9884, 280.02, 279.9637, 280.048, 
    279.99, 280.0644, 280.2057, 280.2654, 280.2337, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.7076, 279.5515, 
    279.9362, 280.2022, 280.1342, 280.0256, 279.9871, 280.05, 280.0066, 
    280.0181, 280.1316, 280.1677, 280.278, 280.4358, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.6312, 280.3207, 279.8989, 
    279.1181, 279.0258, 279.4925, 279.7381, 279.9082, 279.8408, 279.8024, 
    279.9927, 280.0458, 279.9801, 279.9821, 280.0492, 280.1129, 280.2386, 
    278.3331, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.2196, 280.1246, 279.8005, 
    279.1123, 278.8437, 279.1069, 279.6183, 279.5983, 279.8805, 279.7144, 
    279.942, 279.9597, 279.94, 279.8758, 279.9336, 279.9093, 279.9661, 
    280.1106, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.2622, 278.6743, 
    278.7288, 279.31, 279.6081, 279.9091, 279.8698, 279.8611, 279.7872, 
    279.8687, 279.8624, 279.8367, 279.7834, 279.7625, 279.9857, 280.11, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.0947, 278.6002, 
    278.7327, 279.1579, 279.6027, 279.8192, 279.8251, 279.7672, 279.6721, 
    279.7257, 279.7633, 279.7348, 279.7007, 279.7422, 279.9386, 280.0785, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.9955, 278.2114, 
    278.8325, 279.7838, 279.7758, 279.6287, 279.6693, 279.6376, 279.6057, 
    279.6415, 279.6831, 279.7896, 279.781, 279.7464, 279.9234, 280.1089, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.8296, 278.6555, 
    277.7087, 278.5214, 279.7376, 279.6648, 279.1605, 279.1765, 279.1806, 
    279.4865, 279.5964, 279.6723, 279.9641, 279.8994, 279.8259, 280.0058, 
    279.6125, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.9408, 278.4337, 
    278.7756, 279.459, 279.4934, 278.881, 278.5921, 278.9276, 279.3585, 
    279.5063, 279.642, 279.9106, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.3772, _, _, 
    279.7184, 279.6171, 279.3585, 278.8056, 278.6183, 279.017, 279.3239, 
    279.3802, 279.5178, 279.7747, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.3594, 
    279.0207, 278.5473, 278.6123, 279.1168, 279.2466, 279.2576, 279.5351, 
    277.386, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.1797, 
    278.4743, 278.2842, 278.2669, 279.0653, 279.1484, 279.0814, 279.5071, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.1567, 
    278.1678, 277.8053, 278.0629, 278.7706, 278.8426, 279.0135, 279.3784, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 278.4193, 278.416, 278.5337, 278.4522, 278.5168, 
    279.3383, _, _, 279.4039, _, _, 278.2514, 278.1341, 277.798, 277.4796, 
    278.1788, 278.4774, 278.4341, 278.9433, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 278.0911, 278.2601, 278.0482, 278.4938, 278.6233, 
    278.5898, 279.2477, _, _, _, _, _, 278.0863, 277.6967, 277.369, 277.1114, 
    278.2672, 278.8993, 278.7827, 279.085, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 277.774, 277.7, 277.5289, 278.0371, 278.434, 
    278.5336, 278.9521, _, _, _, _, _, 278.5209, 277.9786, 277.2736, 277.084, 
    278.2853, 279.0635, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 277.7354, 277.6465, 277.9712, 278.1647, 
    278.5814, 279.9866, _, 277.9073, 277.5152, 277.8223, 278.3861, 278.4452, 
    278.0108, 277.4971, 277.6643, 278.507, 278.9389, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, 277.9853, 278.4406, 277.9028, 278.6749, _, _, 
    277.8709, 277.2195, 277.4784, 277.6751, 277.5956, 277.5254, 277.4374, 
    277.7198, 278.457, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.9267, _, _, 277.5161, 
    277.2637, 277.2206, 276.7238, 277.2001, 277.3651, 277.6006, 278.3892, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.9645, 278.2161, 277.9534, 
    277.461, 277.3008, 277.3691, 277.2503, 277.1311, 277.3812, 277.9829, 
    278.4565, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 278.1922, _, 277.7226, 277.3818, 
    277.268, 277.2746, 277.4548, 277.5714, 277.5052, 277.757, 276.0721, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.5823, 275.8397, 276.413, 
    276.6071, 277.1882, 277.6274, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.2188, 277.02, 276.0341, 
    274.3827, 274.5943, 275.6299, 276.3824, 276.8616, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 278.8594, 277.4691, 276.8148, 
    275.1505, 273.5242, 273.5737, 274.3829, 275.7479, 276.6379, 276.533, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.8828, 276.2522, 274.3347, 
    273.1601, 273.0244, 273.3189, 274.4734, 275.2237, 275.7833, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.9274, 273.4467, 274.248, 
    273.9681, 273.4105, 272.8058, 273.9072, 275.2976, 276.5013, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.6712, 275.8814, 274.1224, 
    273.9586, 274.538, 274.6036, 274.5869, 274.7482, 275.4168, 276.4592, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 279.3687, _, 277.2096, 276.7476, 276.0802, 
    274.665, 274.0338, 274.8314, 275.4641, 275.6916, 275.8451, 276.0451, 
    276.545, 278.2035, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 276.6808, _, 276.9684, _, 277.1086, 
    275.3448, 274.4252, 274.7439, 275.8261, 276.6003, 277.6399, 276.8841, 
    276.8797, 277.1765, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 277.2939, 277.4904, _, _, 276.7659, 
    276.1925, 274.9077, 274.8026, 276.7263, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 275.6916, 278.5022, _, _, 276.78, 
    275.853, 275.2028, 275.5123, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 276.0755, 277.0032, _, _, 277.1172, 
    275.987, 275.7529, 275.7403, 275.7343, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.6198, 276.266, 
    276.3721, 276.6024, 280.2881, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.8288, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.5026, 
    277.374, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    277.3653, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.5935, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.3125, 275.9853, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.5005, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 278.9684, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.5011, 281.2123, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.7844, 281.1698, 280.8033, 
    280.2764, 280.8499, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.0322, 280.5294, 
    280.3057, 280.722, 280.4402, 280.6487, 280.7616, 280.6664, 280.8568, 
    280.6219, 280.7402, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.9634, 280.6443, 
    280.5098, 280.6756, 280.7571, 280.7148, 280.6152, 280.6536, 280.6294, 
    280.562, 280.5633, 280.4805, 280.4765, 280.5903, 277.5443, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.0678, 280.9941, 
    280.8706, 280.8552, 280.6302, 280.5993, 280.6434, 280.6884, 280.4785, 
    280.5861, 280.5583, 280.6422, 280.7068, 280.6985, 280.6463, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.7471, 
    281.0009, 280.7235, 280.6867, 280.503, 280.5006, 280.4431, 280.5449, 
    280.5213, 280.6361, 280.8422, 280.9159, 280.7782, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.1986, 280.0903, 
    280.4848, 280.7772, 280.6957, 280.5697, 280.4991, 280.5132, 280.4444, 
    280.4677, 280.6133, 280.7012, 280.8574, 281.0151, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.9156, 280.6992, 280.3931, 
    279.6996, 279.5609, 280.0009, 280.2198, 280.4012, 280.3249, 280.2587, 
    280.414, 280.4514, 280.4009, 280.446, 280.5729, 280.6732, 280.7462, 
    279.1562, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.2159, 280.5352, 280.2885, 
    279.6965, 279.3784, 279.5846, 280.0756, 280.0201, 280.2927, 280.1205, 
    280.3473, 280.3579, 280.3552, 280.3395, 280.4621, 280.4844, 280.5182, 
    280.5537, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.7788, 279.2412, 
    279.227, 279.7625, 280.0115, 280.2857, 280.2589, 280.2661, 280.193, 
    280.2849, 280.323, 280.3548, 280.3481, 280.3004, 280.471, 280.5028, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.6616, 279.1917, 
    279.284, 279.6278, 280.011, 280.201, 280.2072, 280.1592, 280.067, 
    280.1321, 280.2088, 280.2351, 280.2424, 280.295, 280.4583, 280.4886, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.5321, 278.821, 
    279.3964, 280.2812, 280.2211, 280.0367, 280.0357, 280.0011, 279.9706, 
    280.0275, 280.1122, 280.2567, 280.2758, 280.2541, 280.4095, 280.4643, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.0455, 279.1322, 
    278.3156, 279.0584, 280.2136, 280.1324, 279.5986, 279.5238, 279.5005, 
    279.8178, 279.95, 280.0564, 280.3588, 280.3508, 280.2482, 280.3563, 
    279.8247, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.3881, 278.9756, 
    279.2557, 279.8975, 279.9382, 279.287, 278.9268, 279.2592, 279.6728, 
    279.8203, 279.9691, 280.2205, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.6189, _, _, 
    280.1237, 279.9874, 279.7458, 279.1209, 278.8993, 279.3155, 279.6158, 
    279.6761, 279.8044, 280.0402, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.616, 
    279.2709, 278.7725, 278.8705, 279.3883, 279.518, 279.53, 279.7495, 
    278.5507, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.3962, 
    278.6471, 278.4622, 278.5004, 279.3355, 279.4171, 279.325, 279.6608, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.6959, 
    278.381, 277.998, 278.3055, 279.0616, 279.1095, 279.2248, 279.5205, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 279.7153, 279.6202, 279.6673, 279.3893, 
    279.2744, 279.8782, _, _, 279.5369, _, _, 278.4398, 278.3774, 278.0803, 
    277.7676, 278.5065, 278.796, 278.7156, 279.1323, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 279.464, 279.59, 279.2377, 279.6232, 279.6057, 
    279.4167, 279.9291, _, _, _, _, _, 278.3509, 278.0164, 277.7704, 
    277.5424, 278.722, 279.2941, 279.0963, 279.2829, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 279.1853, 279.0763, 278.7708, 279.1875, 279.4829, 
    279.4467, 279.7978, _, _, _, _, _, 278.8427, 278.3995, 277.7732, 
    277.6127, 278.8199, 279.5049, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 279.1821, 278.9993, 279.248, 279.3219, 279.6345, 
    280.6498, _, 278.3132, 277.9007, 278.1552, 278.6941, 278.8461, 278.5216, 
    278.0922, 278.2733, 279.0472, 279.421, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, 279.4219, 279.8371, 279.1386, 279.832, _, _, 
    278.4427, 277.7812, 278.0182, 278.1919, 278.1286, 278.1567, 278.133, 
    278.4279, 279.078, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.6852, _, _, 278.2364, 
    277.9868, 277.9293, 277.4465, 278.0132, 278.1859, 278.4128, 279.1088, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.922, 279.0373, 278.8334, 
    278.3731, 278.1604, 278.2397, 278.1636, 278.1003, 278.3551, 278.8667, 
    279.2491, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 279.1503, _, 278.6428, 278.3754, 
    278.2881, 278.2707, 278.4546, 278.5892, 278.5212, 278.7388, 276.2067, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.657, 277.0777, 277.6246, 
    277.7661, 278.2868, 278.6543, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.14, 278.0123, 277.2431, 
    275.8255, 276.0841, 276.9782, 277.5993, 278.0031, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 279.8585, 278.5143, 277.8541, 
    276.6003, 275.3235, 275.3702, 276.0347, 277.1447, 277.8805, 278.1903, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.9865, 277.4166, 275.7661, 
    274.4071, 274.6668, 275.1909, 275.9403, 276.6217, 277.0569, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.9984, 274.8752, 275.8742, 
    275.6248, 275.2773, 273.9154, 275.4643, 276.6918, 277.7506, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.7697, 277.1775, 275.767, 
    275.6852, 276.3089, 276.3977, 276.3395, 276.363, 276.9024, 277.8336, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 279.9155, _, 278.4607, 277.9834, 277.4978, 
    276.3113, 275.7999, 276.7405, 277.4366, 277.5555, 277.5366, 277.6123, 
    278.011, 279.1763, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 277.9758, _, 278.2606, _, 278.3976, 
    277.0487, 276.2654, 276.652, 277.8276, 278.6102, 278.7449, 278.783, 
    278.3453, 278.1653, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 278.5714, 278.6169, _, _, 277.9743, 
    277.8506, 276.6547, 276.6455, 278.2296, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 277.5676, 278.7439, _, _, 278.0752, 
    277.5104, 276.971, 277.3331, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 277.7649, 278.3937, _, _, 278.5212, 
    277.4829, 277.3661, 277.4718, 277.4604, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.6383, 277.8439, 
    278.0234, 278.271, 280.7772, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.3543, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.5524, 
    278.5982, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    278.4551, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    277.0438, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.6083, 275.9683, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.0872, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 277.8929, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.0008, 279.7851, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.5722, 279.5775, 279.1222, 
    278.4014, 279.2239, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.4051, 278.7635, 
    278.4308, 278.9356, 278.8593, 278.7015, 278.7767, 278.7241, 279.6156, 
    278.7227, 278.9314, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.1434, 278.6037, 
    278.4619, 278.6759, 278.7415, 278.669, 278.5629, 278.6536, 278.6818, 
    278.6169, 278.7089, 278.7132, 278.7932, 279.028, 276.4333, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.008, 278.9279, 
    278.7455, 278.7068, 278.4778, 278.3802, 278.3752, 278.4162, 278.3611, 
    278.6248, 278.7101, 278.8984, 279.1108, 279.3264, 279.5475, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.9024, 
    278.7607, 278.4762, 278.4095, 278.1539, 278.25, 278.4174, 278.7091, 
    278.8045, 279.0149, 279.2969, 279.4778, 279.5732, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.7041, 278.1278, 
    278.4145, 278.7018, 278.6086, 278.4616, 278.4174, 278.5652, 278.6541, 
    278.8033, 279.0369, 279.1985, 279.4152, 279.6453, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.5633, 279.3366, 278.8042, 
    277.8665, 277.5996, 278.0172, 278.2366, 278.4615, 278.442, 278.4449, 
    278.7003, 278.8113, 278.8222, 278.9249, 279.0907, 279.2327, 279.4291, 
    278.2753, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.8812, 279.1046, 278.5801, 
    277.7873, 277.3502, 277.5003, 278.0866, 278.1305, 278.5193, 278.3985, 
    278.6933, 278.7671, 278.7867, 278.7785, 278.9286, 278.9593, 279.0416, 
    279.2321, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.8328, 277.1678, 
    277.1437, 277.7779, 278.1678, 278.5582, 278.5612, 278.6147, 278.5949, 
    278.7013, 278.7275, 278.7493, 278.7401, 278.6887, 278.9296, 279.0871, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.5793, 277.0639, 
    277.1583, 277.6107, 278.2014, 278.5158, 278.5667, 278.5465, 278.4626, 
    278.5204, 278.5628, 278.5459, 278.5519, 278.6058, 278.7989, 278.9557, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.528, 276.7139, 
    277.3174, 278.3903, 278.4873, 278.4328, 278.5064, 278.4696, 278.3941, 
    278.4048, 278.4391, 278.5645, 278.5757, 278.5319, 278.6707, 278.877, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.5373, 277.2818, 
    276.264, 277.0303, 278.4069, 278.4821, 278.0999, 278.1065, 278.0564, 
    278.3036, 278.3762, 278.4406, 278.7303, 278.6794, 278.5869, 278.741, 
    278.4312, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.5681, 277.0318, 
    277.3946, 278.2012, 278.4077, 277.8766, 277.5004, 277.795, 278.2024, 
    278.3282, 278.4366, 278.6635, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.2768, _, _, 
    278.4483, 278.5028, 278.4215, 277.8428, 277.5253, 277.8772, 278.1903, 
    278.2429, 278.3364, 278.5466, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.3636, 
    278.2363, 277.6441, 277.6078, 278.0589, 278.1907, 278.1772, 278.3805, 
    277.1379, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.3466, 
    277.7388, 277.4542, 277.3726, 278.1203, 278.1942, 278.0535, 278.3705, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.5154, 
    277.4668, 277.0136, 277.1962, 277.8877, 277.9103, 277.9748, 278.2583, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 278.6624, 278.4802, 278.3907, 278.0195, 
    278.0018, 279.0532, _, _, 278.6561, _, _, 277.5242, 277.5072, 277.1349, 
    276.654, 277.2859, 277.516, 277.3915, 277.8261, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 278.591, 278.6155, 278.2188, 278.5404, 278.4583, 
    278.2767, 279.0847, _, _, _, _, _, 277.2773, 276.9446, 276.6794, 
    276.2112, 277.3354, 277.8332, 277.6064, 277.853, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 278.4282, 278.2177, 277.8536, 278.2445, 278.5188, 
    278.4816, 278.9269, _, _, _, _, _, 277.8209, 277.2644, 276.5096, 
    276.0852, 277.2503, 277.9766, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 278.3532, 278.0749, 278.2958, 278.3917, 
    278.7705, 279.2757, _, 277.1288, 276.959, 277.3228, 277.7871, 277.928, 
    277.4147, 276.7513, 276.7397, 277.4897, 277.8994, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, 278.4986, 278.9029, 278.2445, 279.0162, _, _, 
    277.4317, 276.8596, 277.1039, 277.2438, 277.117, 276.9282, 276.735, 
    276.9187, 277.5545, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.3164, _, _, 277.2761, 
    276.9854, 276.8325, 276.1796, 276.6447, 276.7362, 276.863, 277.5983, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.4241, 278.1666, 278.0707, 
    277.5483, 277.1992, 277.113, 276.8257, 276.675, 276.8795, 277.3551, 
    277.7678, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 278.6197, _, 277.9774, 277.7389, 
    277.5739, 277.4077, 277.4036, 277.3419, 277.1003, 277.2514, 275.5806, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.1197, 276.7209, 277.0714, 
    276.9524, 277.2912, 277.4909, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.6452, 277.6425, 276.9257, 
    275.4874, 275.462, 276.0885, 276.546, 276.8085, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 279.0268, 277.2972, 277.6117, 
    276.2909, 274.7977, 274.7185, 275.1063, 276.057, 276.82, 276.3434, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.87, 277.303, 275.5406, 
    274.2962, 274.1021, 274.2278, 274.9091, 275.3836, 275.6811, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.6466, 274.7459, 275.3047, 
    274.8152, 274.2241, 273.2891, 273.9655, 275.0133, 276.114, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.3401, 277.0669, 275.5009, 
    275.074, 275.3581, 275.1324, 274.8372, 274.6754, 275.1092, 276.0621, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 278.0139, _, 276.8508, 277.7931, 277.3652, 
    276.0366, 275.2156, 275.666, 275.9924, 275.8892, 275.6456, 275.7188, 
    276.2417, 279.1501, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 277.7852, _, 277.837, _, 276.8471, 
    276.5578, 275.5607, 275.5967, 276.4659, 276.9769, 278.1729, 277.0541, 
    276.6372, 276.9848, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 277.1519, 278.136, _, _, 278.1725, 
    277.179, 275.8249, 275.5336, 277.1818, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 276.3171, 277.8159, _, _, 277.5974, 
    276.638, 275.8526, 276.0417, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 276.4314, 277.8945, _, _, 278.152, 
    276.507, 276.2739, 276.2951, 276.2446, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.7834, 276.6893, 
    276.9337, 277.2144, 278.7738, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.3549, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.6879, 
    277.2361, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    277.6372, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.5223, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.0873, 275.3484, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.1738, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 284.4954, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.9373, 285.0029, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.4349, 285.3036, 285.2369, 
    284.6889, 285.3124, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.208, 284.8527, 
    284.6528, 285.3537, 284.696, 286.397, 286.0988, 286.2746, 285.7757, 
    285.6713, 286.0729, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.2647, 285.0791, 
    285.1833, 285.7264, 286.1018, 286.1677, 286.1681, 286.3518, 286.2937, 
    286.0111, 286.0122, 285.9332, 285.882, 285.8437, 283.6741, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.4755, 285.5856, 
    285.8462, 286.1399, 286.0662, 286.0663, 286.1774, 286.2653, 285.8317, 
    285.8468, 285.6821, 285.7336, 285.6586, 285.5551, 285.2408, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.0386, 
    286.2914, 286.1531, 286.1722, 285.9246, 285.9163, 285.7319, 285.7026, 
    285.4729, 285.4727, 285.5918, 285.4424, 285.0423, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.0782, 285.4648, 
    285.7542, 286.1786, 286.1809, 286.0554, 285.955, 285.9366, 285.7163, 
    285.567, 285.6129, 285.5681, 285.6371, 285.6759, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.9034, 285.9152, 285.8654, 
    285.0992, 284.895, 285.3648, 285.6308, 285.9058, 285.8093, 285.7104, 
    285.8297, 285.7146, 285.4792, 285.3988, 285.4491, 285.4772, 285.4636, 
    284.6622, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.8377, 285.6003, 285.4849, 
    284.9834, 284.6436, 284.8702, 285.4771, 285.4504, 285.8213, 285.5611, 
    285.7082, 285.5442, 285.3755, 285.2052, 285.288, 285.2602, 285.2686, 
    285.1245, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.9368, 284.4414, 
    284.4302, 285.0971, 285.4469, 285.802, 285.6976, 285.5608, 285.2905, 
    285.2422, 285.1492, 285.1223, 285.0885, 284.9897, 285.0578, 284.9126, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.9388, 284.3872, 
    284.4521, 284.848, 285.3605, 285.6252, 285.5872, 285.3862, 285.1024, 
    285.0139, 284.9646, 284.9388, 284.9296, 284.9345, 285.0109, 284.9017, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.0005, 284.065, 
    284.5863, 285.551, 285.5115, 285.3965, 285.4022, 285.2119, 285.0029, 
    284.8695, 284.8113, 284.9033, 284.8734, 284.8026, 284.8637, 284.7851, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.7232, 284.6953, 
    283.591, 284.2607, 285.5286, 285.4268, 284.9052, 284.907, 284.702, 
    284.8862, 284.8429, 284.7246, 284.8985, 284.875, 284.6708, 284.657, 
    284.3421, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.8831, 284.3129, 
    284.5346, 285.2147, 285.288, 284.6066, 284.19, 284.4175, 284.7759, 
    284.8028, 284.6891, 284.5961, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.9476, _, _, 
    285.4174, 285.3182, 285.1773, 284.5271, 284.1888, 284.5338, 284.7806, 
    284.6547, 284.4321, 284.3849, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.1336, 
    284.824, 284.2979, 284.2684, 284.7192, 284.7193, 284.4857, 284.3696, 
    283.092, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.9718, 
    284.339, 284.1224, 283.9718, 284.6892, 284.6166, 284.24, 284.3203, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.8764, 
    284.1927, 283.6906, 283.7867, 284.3639, 284.2141, 284.0622, 284.204, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 284.5874, 284.6594, 284.8378, 284.6763, 
    284.5812, 285.2396, _, _, 284.8876, _, _, 284.6142, 284.4153, 283.9829, 
    283.4426, 283.947, 283.9872, 283.6091, 283.7654, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 284.216, 284.5397, 284.2917, 284.9924, 285.1198, 
    284.8754, 285.2724, _, _, _, _, _, 284.4025, 283.9417, 283.7213, 
    283.1382, 283.9642, 284.2089, 283.653, 283.6337, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 283.9789, 284.0299, 283.868, 284.5545, 284.9985, 
    284.8667, 285.1087, _, _, _, _, _, 284.877, 284.3718, 283.6673, 283.085, 
    283.788, 284.1305, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 284.2325, 284.162, 284.5922, 284.7034, 284.9211, 
    285.7315, _, 284.2892, 283.9397, 284.2292, 284.8193, 285.0197, 284.6009, 
    283.946, 283.6272, 283.7878, 283.8586, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, 284.3773, 284.9957, 284.2049, 284.8137, _, _, 
    284.3432, 283.868, 284.2329, 284.4677, 284.353, 284.2864, 283.9503, 
    283.6407, 283.5834, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.0387, _, _, 284.3932, 
    284.2941, 284.2758, 283.5501, 284.1002, 283.9196, 283.4344, 283.4143, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.8069, 284.688, 284.8562, 
    284.6363, 284.5474, 284.6624, 284.4498, 284.073, 283.8209, 283.6728, 
    283.467, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 284.1845, _, 284.4485, 284.4078, 
    284.589, 284.6484, 284.7991, 284.7875, 284.245, 283.8524, 280.0029, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.8759, 283.4433, 284.1074, 
    284.0847, 284.4531, 284.5127, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.0209, 283.9028, 283.5666, 
    282.4197, 282.6277, 283.2371, 283.556, 283.449, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 285.102, 283.542, 283.7624, 
    283.0285, 282.0125, 282.0339, 282.3698, 283.1276, 283.4125, 284.3994, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.9919, 283.4377, 282.4964, 
    281.7614, 281.7885, 281.8981, 282.3833, 282.5479, 282.3879, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.8368, 281.9449, 283.1948, 
    283.007, 282.4922, 281.4861, 281.8282, 282.4912, 282.8781, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.3747, 283.2695, 282.6701, 
    282.9024, 283.7654, 283.828, 283.5661, 283.111, 283.0041, 283.2098, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 285.4368, _, 283.2258, 283.4045, 283.5949, 
    283.1272, 282.8841, 284.0382, 284.8403, 284.8476, 284.4295, 283.8287, 
    283.5258, 283.2982, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 283.4608, _, 283.2983, _, 283.2421, 
    283.5634, 283.2005, 283.4805, 284.8892, 285.6749, 283.2839, 285.3781, 
    283.8532, 282.8722, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 283.4695, 283.2341, _, _, 283.0997, 
    284.045, 283.1132, 283.0863, 283.4499, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 284.1464, 284.563, _, _, 282.9432, 
    283.696, 283.3829, 283.7865, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 283.9155, 283.2917, _, _, 283.4019, 
    283.476, 283.5676, 283.7939, 283.4847, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.9722, 283.3239, 
    284.255, 284.1536, 286.0193, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.6312, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.186, 
    283.3353, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    283.0565, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    281.9973, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    281.3661, 280.0912, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.7614, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 285.5234, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.0261, 287.162, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.6175, 287.5185, 287.8371, 
    287.5563, 288.3271, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.1142, 287.1256, 
    287.4058, 288.2428, 289.4631, 289.2658, 288.7545, 288.9729, 286.8089, 
    288.2659, 289.6769, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.2204, 287.4623, 
    287.7634, 288.2206, 288.595, 288.7958, 288.9529, 289.3281, 289.5509, 
    289.6589, 289.991, 290.2057, 290.4017, 290.631, 283.0873, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.4618, 287.8947, 
    288.2582, 288.6066, 288.6617, 288.931, 289.3121, 289.6907, 289.6806, 
    290.037, 290.2041, 290.5128, 290.6465, 290.6428, 290.3186, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.5452, 
    288.7569, 288.7105, 289.0221, 289.171, 289.5578, 289.765, 290.0876, 
    290.2041, 290.4913, 290.782, 290.7374, 290.344, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.1566, 287.3222, 
    287.9651, 288.6482, 288.7683, 288.8872, 289.1914, 289.5946, 289.8174, 
    290.0574, 290.4212, 290.6888, 290.8913, 290.9468, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.0042, 286.9716, 287.0056, 
    286.5533, 286.8167, 287.7013, 288.1765, 288.5648, 288.6834, 288.9466, 
    289.4898, 289.8111, 289.9481, 290.1873, 290.4953, 290.6779, 290.6842, 
    285.4996, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.8047, 286.4621, 286.5428, 
    286.518, 286.6836, 287.3509, 288.1993, 288.2499, 288.7813, 288.7627, 
    289.3293, 289.5938, 289.7666, 289.9013, 290.2001, 290.3228, 290.401, 
    290.2444, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.337, 286.4194, 
    286.869, 287.8532, 288.367, 288.8816, 288.939, 289.0923, 289.2356, 
    289.5438, 289.7238, 289.8649, 289.9667, 289.9909, 290.2166, 289.9934, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.3854, 286.2713, 
    286.8865, 287.6189, 288.3679, 288.8098, 288.8994, 288.893, 288.9245, 
    289.1826, 289.4036, 289.491, 289.5908, 289.8042, 290.0945, 289.9785, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.1814, 285.8199, 
    287.0498, 288.4112, 288.5112, 288.5608, 288.754, 288.7378, 288.7267, 
    288.8743, 289.0174, 289.2084, 289.285, 289.4099, 289.7212, 289.6857, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.2846, 285.6412, 
    285.1439, 286.5637, 288.315, 288.2611, 287.8782, 288.1484, 288.201, 
    288.5337, 288.7, 288.7691, 288.9678, 289.1501, 289.0573, 289.1915, 
    287.8334, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.7727, 285.7673, 
    286.5767, 287.6432, 287.8878, 287.3711, 287.25, 287.8294, 288.346, 
    288.4512, 288.5155, 288.563, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.719, _, _, 287.2391, 
    287.3734, 287.4522, 287.0206, 287.0723, 287.7908, 288.1985, 288.1301, 
    288.0313, 288.1595, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.684, 
    286.653, 286.432, 286.9434, 287.7627, 287.9847, 287.8632, 287.8031, 
    285.45, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.1821, 
    285.7337, 286.0001, 286.366, 287.5529, 287.7562, 287.5398, 287.6409, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.0822, 
    285.3294, 285.3325, 286.0008, 287.0475, 287.1992, 287.2733, 287.4689, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 286.2361, 286.3193, 286.4856, 286.2663, 
    286.1336, 286.7625, _, _, 285.9271, _, _, 285.0929, 285.0836, 284.9547, 
    284.9731, 286.1063, 286.5003, 286.4513, 286.9591, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 285.5769, 285.938, 285.7474, 286.4272, 286.523, 
    286.3137, 286.7457, _, _, _, _, _, 284.9459, 284.6198, 284.6608, 
    284.6976, 286.207, 286.847, 286.575, 286.9051, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, 285.0445, 285.1225, 285.0196, 285.7481, 286.2202, 
    286.1667, 286.4598, _, _, _, _, _, 285.583, 285.1486, 284.6732, 284.6704, 
    286.1768, 286.8997, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 284.9945, 284.9694, 285.4403, 285.6932, 286.077, 
    290.687, _, 285.3647, 284.971, 285.212, 285.6855, 285.7846, 285.389, 
    285.0649, 285.4486, 286.3152, 286.6804, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, 284.8777, 285.5258, 285.0264, 285.8229, _, _, 
    285.2335, 284.8015, 285.2351, 285.3577, 285.1586, 285.0504, 285.1145, 
    285.5691, 286.2523, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.2716, _, _, 285.3337, 
    285.2601, 285.1444, 284.4141, 285.0305, 285.2496, 285.4355, 286.1943, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.0013, 285.6929, 285.9662, 
    285.634, 285.495, 285.5718, 285.338, 285.1425, 285.4315, 285.9576, 
    286.2501, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 284.7314, _, 285.3206, 285.4491, 
    285.6112, 285.6514, 285.8399, 285.8736, 285.5601, 285.7333, 282.0126, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.306, 284.1358, 284.971, 
    285.1119, 285.6373, 285.8607, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.1079, 284.0836, 283.7308, 
    282.9565, 283.4535, 284.326, 284.871, 285.1314, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 286.3276, 285.6212, 283.7508, 
    283.1139, 282.3795, 282.7501, 283.4583, 284.6308, 285.3387, 285.3276, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.2069, 283.2269, 282.4953, 
    281.9975, 282.24, 282.7087, 283.7133, 284.1986, 284.3841, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.3146, 281.852, 283.1808, 
    283.04, 282.8222, 282.3705, 283.1411, 284.3355, 285.2567, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.9758, 283.1267, 282.3441, 
    282.7135, 283.6832, 283.8772, 284.0004, 284.0992, 284.5805, 285.3595, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 286.9834, _, 285.7414, 283.3557, 283.2821, 
    282.6563, 282.5381, 283.9793, 284.9102, 285.0236, 284.9848, 284.9786, 
    285.309, 283.9461, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 283.3578, _, 283.4039, _, 285.4762, 
    282.9262, 282.7375, 283.47, 285.1009, 285.8674, 283.6351, 285.813, 
    285.4479, 285.4137, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 285.4304, 283.5518, _, _, 283.2774, 
    283.412, 282.6978, 283.0675, 284.1529, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 284.3936, 285.5286, _, _, 283.0332, 
    283.1826, 283.1156, 283.8129, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 284.2635, 283.4037, _, _, 283.5495, 
    282.9497, 283.0663, 283.509, 283.6461, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.8396, 283.9873, 
    283.8456, 284.1613, 288.6338, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.1205, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.809, 
    285.4108, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    283.6279, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    282.5311, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    282.2342, 281.8941, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 294.1141, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 289.1718, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.7405, 292.1293, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 296.0645, 292.841, 293.7014, 
    293.9014, 294.0972, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.3386, 292.7533, 
    293.2753, 294.2085, 293.9911, 297, 295.8654, 296.4326, 291.8285, 
    294.6871, 297.0214, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.5709, 293.2369, 
    293.8943, 294.7183, 295.523, 296.0438, 296.4758, 297.0791, 297.4254, 
    297.4051, 297.6319, 297.9148, 298.227, 298.4543, 285.9212, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 293.0215, 293.7612, 
    294.7737, 295.5681, 296.0978, 296.5531, 297.0514, 297.4786, 297.5029, 
    297.7983, 297.8997, 298.1832, 298.2755, 298.0072, 296.8398, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 296.9357, 
    295.8319, 296.3208, 296.7845, 296.9977, 297.311, 297.4712, 297.7395, 
    297.7917, 297.9005, 298.0209, 297.6272, 296.291, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.1727, 294.2439, 
    294.9181, 295.949, 296.4442, 296.7588, 297.0359, 297.307, 297.4104, 
    297.5435, 297.7596, 297.7952, 297.6982, 297.3226, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.0975, 292.5047, 293.1029, 
    293.1248, 293.6868, 294.8661, 295.7139, 296.3542, 296.6233, 296.8168, 
    297.1858, 297.3778, 297.3911, 297.4424, 297.5069, 297.3457, 296.6568, 
    289.1045, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.4341, 291.8948, 292.455, 
    292.8079, 293.3619, 294.4461, 295.6105, 295.9551, 296.6236, 296.6331, 
    297.0246, 297.2024, 297.2801, 297.2214, 297.2685, 297.0719, 296.5823, 
    295.3923, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.2513, 293.0027, 
    293.9046, 295.1262, 295.8319, 296.4765, 296.6418, 296.7775, 296.8863, 
    297.1287, 297.1359, 297.0366, 296.8148, 296.273, 295.7518, 294.6631, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.707, 292.8905, 
    293.744, 294.6592, 295.5553, 296.1288, 296.3815, 296.504, 296.6032, 
    296.8579, 296.9478, 296.7919, 296.5078, 296.1347, 295.6856, 294.7282, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.6748, 292.4643, 
    293.7119, 295.1377, 295.391, 295.6512, 296.0075, 296.2093, 296.3681, 
    296.5771, 296.6631, 296.5345, 296.135, 295.6731, 295.259, 294.2902, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.7337, 291.9539, 
    291.6102, 292.9659, 294.7182, 294.8687, 294.8406, 295.2299, 295.4819, 
    296.0465, 296.2851, 296.2218, 295.9561, 295.8504, 295.0689, 294.3624, 
    293.8385, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.7473, 291.7265, 
    292.5043, 293.6861, 294.2818, 294.2126, 294.3438, 294.9388, 295.628, 
    295.8258, 295.6086, 294.9414, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.315, _, _, 292.5554, 
    293.1086, 293.7615, 293.8197, 294.0544, 294.7427, 295.2452, 295.2226, 
    294.7089, 294.2633, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.5549, 
    293.1364, 293.293, 293.8065, 294.5671, 294.8315, 294.6096, 293.9038, 
    288.1628, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.9, 
    292.403, 292.8521, 293.1447, 294.2411, 294.425, 293.9263, 293.2617, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 294.9114, 
    292.0917, 292.1966, 292.8001, 293.7199, 293.7248, 293.2802, 292.8942, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 289.9971, 290.2084, 290.464, 290.3806, 290.262, 
    290.4582, _, _, 290.2698, _, _, 291.5617, 291.7162, 291.7819, 291.7904, 
    292.7546, 293.0631, 292.7872, 292.5838, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 289.1241, 289.6299, 289.5406, 290.2859, 290.4388, 
    290.1599, 290.3153, _, _, _, _, _, 291.3478, 291.2292, 291.4124, 291.268, 
    292.5233, 292.9964, 292.3649, 292.0424, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 288.5088, 288.725, 288.7047, 289.4595, 289.895, 
    289.7409, 289.9081, _, _, _, _, _, 291.7491, 291.5871, 291.2158, 
    290.9133, 291.9197, 292.4393, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 288.4765, 288.4728, 288.9344, 289.0941, 
    289.3337, 298.2717, _, 290.0002, 289.9064, 290.5951, 291.4253, 291.9028, 
    291.7639, 291.377, 291.3066, 291.6131, 291.7356, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, 288.0456, 288.6103, 288.0633, 288.6244, _, _, 
    289.4816, 289.4513, 290.4388, 291.0482, 291.2435, 291.3737, 291.3202, 
    291.2579, 291.1993, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.4916, _, _, 289.7179, 
    290.1654, 290.5652, 290.2842, 291.0979, 291.237, 290.9697, 290.9062, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.8255, 289.3395, 289.8391, 
    289.8842, 290.154, 290.6661, 290.8286, 290.8423, 290.9618, 291.0188, 
    290.7881, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 288.0262, _, 288.9574, 289.29, 
    289.8169, 290.1773, 290.6635, 290.953, 290.7686, 290.686, 283.4617, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.1447, 288.1986, 289.372, 
    289.6873, 290.3685, 290.6349, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.6543, 287.8914, 287.6059, 
    287.0405, 287.8491, 288.8976, 289.5415, 289.7145, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 289.5497, 289.9067, 287.4436, 
    287.0089, 286.4873, 287.0969, 287.8788, 289.0047, 289.6267, 288.385, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.4324, 286.6989, 286.3912, 
    286.1417, 286.5554, 287.0741, 288.0075, 288.4554, 288.5005, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.075, 285.7678, 287.5537, 
    287.4701, 287.1799, 286.5703, 287.2608, 288.1619, 288.7078, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.0437, 286.3915, 286.2955, 
    286.9061, 287.9366, 288.0459, 288.0058, 287.8738, 288.0336, 288.4706, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 294.0276, _, 288.6398, 286.2251, 286.5561, 
    286.4562, 286.5344, 287.8948, 288.7418, 288.7762, 288.5534, 288.2137, 
    288.2289, 286.2427, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 286.2591, _, 286.0636, _, 288.2309, 
    286.5208, 286.548, 287.1331, 288.5672, 289.126, 286.1544, 288.7925, 
    288.2361, 289.3455, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 288.0631, 286.1037, _, _, 286.0705, 
    286.7701, 286.1187, 286.4915, 286.6264, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 287.6348, 292.084, _, _, 285.6241, 
    286.3089, 286.342, 287.0012, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 287.3455, 285.9029, _, _, 285.9915, 
    285.7983, 286.0106, 286.4978, 286.5739, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.7281, 286.6734, 
    286.6324, 286.7829, 295.5705, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.5397, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.8782, 
    288.036, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    285.6772, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    284.7975, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    284.313, 283.5242, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.9074, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 289.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.7653, 290.8331, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 295.3229, 291.1286, 291.5419, 
    291.6682, 292.3105, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.6721, 290.7755, 
    291.1761, 292.0977, 293.7359, 293.6813, 293.0569, 293.3725, 290.2906, 
    292.3684, 293.8005, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.8335, 291.191, 
    291.6996, 292.3596, 292.8741, 293.1529, 293.353, 293.7292, 293.9813, 
    294.1157, 294.4926, 294.8342, 295.2872, 295.7586, 287.0718, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.1828, 291.7053, 
    292.3872, 292.8897, 293.1376, 293.4011, 293.7421, 294.1034, 294.257, 
    294.6992, 294.9316, 295.4146, 295.7578, 295.8301, 295.1224, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 293.6531, 
    293.0833, 293.3269, 293.6393, 293.7574, 294.0181, 294.2849, 294.7261, 
    294.9312, 295.2802, 295.7681, 295.8463, 295.176, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.7754, 291.5751, 
    292.2823, 293.1365, 293.4541, 293.652, 293.8777, 294.1376, 294.3131, 
    294.6277, 295.065, 295.3959, 295.7245, 295.8348, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.5517, 290.7848, 290.9957, 
    290.7641, 291.1833, 292.1996, 292.8914, 293.3821, 293.5524, 293.7424, 
    294.1396, 294.3682, 294.5401, 294.8485, 295.2237, 295.4859, 295.4829, 
    288.9427, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.9645, 290.3236, 290.5833, 
    290.7206, 291.041, 291.8657, 292.8564, 293.0831, 293.6167, 293.6027, 
    294.0924, 294.2599, 294.4374, 294.6349, 294.9984, 295.1709, 295.2831, 
    294.877, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.4465, 290.7485, 
    291.4052, 292.4754, 293.096, 293.6282, 293.767, 293.9593, 294.0442, 
    294.3156, 294.5368, 294.7464, 294.8509, 294.7861, 294.9298, 294.3999, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.6458, 290.6394, 
    291.369, 292.2294, 293.0253, 293.4884, 293.683, 293.7996, 293.8508, 
    294.0774, 294.2933, 294.3967, 294.4658, 294.5763, 294.7359, 294.383, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.6517, 290.2839, 
    291.4846, 292.9158, 293.1334, 293.282, 293.486, 293.5721, 293.6424, 
    293.7805, 293.9352, 294.0474, 294.0475, 294.0652, 294.2729, 294.0124, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.6052, 290.2473, 
    289.7418, 291.0508, 292.8352, 292.9516, 292.7898, 292.9664, 292.9836, 
    293.359, 293.4989, 293.5284, 293.5585, 293.8047, 293.5055, 293.4883, 
    292.2115, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.3754, 290.3185, 
    291.0401, 292.1578, 292.6355, 292.3617, 292.2053, 292.5768, 293.0595, 
    293.1786, 293.1372, 292.9024, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.679, _, _, 291.4817, 
    291.857, 292.2765, 292.062, 292.0078, 292.4999, 292.8362, 292.8054, 
    292.5718, 292.4272, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291.3429, 
    291.618, 291.5633, 291.8866, 292.4799, 292.5931, 292.4879, 292.2358, 
    287.9111, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.8456, 
    290.7709, 291.0993, 291.3661, 292.3412, 292.4207, 292.1314, 291.9952, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 292.3088, 
    290.3855, 290.3997, 291.0234, 291.9298, 291.9974, 291.8499, 291.8082, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 289.1621, 289.2466, 289.4198, 289.3099, 
    289.2754, 289.7331, _, _, 289.7783, _, _, 290.1388, 290.073, 290.037, 
    290.0007, 290.9585, 291.3488, 291.2468, 291.4022, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 288.6538, 289.0065, 288.7953, 289.4116, 289.5637, 
    289.3871, 289.7088, _, _, _, _, _, 289.9905, 289.6799, 289.76, 289.6047, 
    290.8349, 291.4151, 290.9799, 290.975, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 288.2974, 288.4046, 288.2951, 288.9048, 289.2852, 
    289.1893, 289.4474, _, _, _, _, _, 290.3335, 290.0728, 289.6308, 
    289.4147, 290.5822, 291.2087, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 288.4191, 288.4096, 288.7827, 288.8664, 
    289.1044, 295.8835, _, 289.3907, 288.895, 289.2585, 290.0176, 290.3433, 
    290.1165, 289.7378, 289.8937, 290.5358, 290.8243, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, 288.382, 288.917, 288.276, 288.8513, _, _, 
    289.0302, 288.4583, 289.0679, 289.4957, 289.6044, 289.5726, 289.5298, 
    289.7878, 290.2602, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.4315, _, _, 288.8284, 
    288.8828, 289.0397, 288.6086, 289.247, 289.3531, 289.3863, 289.9735, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.225, 289.0702, 289.22, 
    288.9104, 288.8611, 289.1044, 289.0886, 288.9626, 289.1297, 289.511, 
    289.692, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 288.287, _, 288.6635, 288.6563, 
    288.7645, 288.8137, 289.0484, 289.1607, 288.9265, 288.9978, 284.2264, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.069, 287.5948, 288.2911, 
    288.3784, 288.7779, 288.8703, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.1085, 288.2348, 287.7429, 
    286.6398, 287.0501, 287.7892, 288.1541, 288.1819, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 289.3069, 288.4733, 287.9445, 
    287.201, 286.2769, 286.5225, 287.0288, 287.8932, 288.3923, 288.0266, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.2805, 287.593, 286.6581, 
    286.0097, 286.1366, 286.4639, 287.1237, 287.4077, 287.4701, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.1883, 286.0087, 287.2983, 
    287.0095, 286.6851, 286.0521, 286.4058, 287.2366, 287.9484, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.5754, 287.4589, 286.675, 
    286.8547, 287.5818, 287.5956, 287.5112, 287.276, 287.3912, 287.9368, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 291.2314, _, 288.1901, 287.4968, 287.6488, 
    287.0473, 286.6968, 287.7243, 288.3969, 288.3671, 288.0645, 287.7421, 
    287.8327, 287.155, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 287.5063, _, 287.1884, _, 287.9152, 
    287.3116, 286.9215, 287.1935, 288.37, 288.8617, 287.3599, 288.5733, 
    287.9107, 288.4136, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 287.8205, 287.2887, _, _, 287.0477, 
    287.7599, 286.8296, 286.875, 287.1157, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 287.6453, 290.5301, _, _, 286.8657, 
    287.2977, 287.0471, 287.3091, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 287.3496, 286.9622, _, _, 286.9484, 
    287.0147, 287.0565, 287.2207, 287.0059, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.6078, 287.0047, 
    287.5386, 287.5108, 292.8891, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.1818, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.7697, 
    287.8067, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    286.6235, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    285.6334, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    285.1101, 284.3122, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.8927, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 286.2799, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.9907, 288.7847, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 290.7077, 288.8628, 288.7497, 
    288.3524, 288.7487, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.7689, 288.4397, 
    288.2899, 288.7094, 290.1369, 289.7293, 289.4843, 289.6035, 288.7423, 
    288.7856, 290.0081, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.9061, 288.654, 
    288.5815, 288.9159, 289.3822, 289.6271, 289.6491, 289.7988, 289.9166, 
    289.9549, 290.1162, 290.2507, 290.4729, 290.7428, 285.4664, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.1044, 289.1094, 
    289.1807, 289.5329, 289.6071, 289.7769, 289.9096, 290.087, 289.9878, 
    290.2277, 290.402, 290.7797, 290.8766, 290.8846, 290.7549, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.9453, 
    289.6083, 289.7089, 289.9597, 289.943, 290.0629, 290.0682, 290.2887, 
    290.4329, 290.7807, 291.068, 291.021, 290.7648, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.7879, 288.4102, 
    288.8177, 289.3837, 289.6486, 289.8499, 290.0341, 290.1837, 290.1729, 
    290.2821, 290.5994, 290.8536, 291.056, 291.1166, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.7977, 288.7484, 288.551, 
    288.0717, 288.0376, 288.5955, 289.0372, 289.4903, 289.6938, 289.8456, 
    290.1432, 290.2522, 290.2598, 290.4042, 290.6317, 290.7566, 290.7462, 
    286.3831, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.7065, 288.5864, 288.4673, 
    288.1534, 288.0059, 288.3872, 289.0408, 289.2196, 289.7986, 289.7832, 
    290.1183, 290.1845, 290.237, 290.2665, 290.4449, 290.4846, 290.4336, 
    290.2262, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.1939, 287.8876, 
    288.1086, 288.8486, 289.3406, 289.8513, 289.9823, 290.0826, 290.0439, 
    290.1831, 290.2519, 290.3052, 290.2923, 290.1172, 290.1813, 290.0716, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.1877, 287.8539, 
    288.1921, 288.7621, 289.3764, 289.796, 289.9995, 290.06, 289.9755, 
    290.0363, 290.1213, 290.135, 290.1301, 290.141, 290.2188, 290.1391, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.0773, 287.5098, 
    288.339, 289.4644, 289.5454, 289.6399, 289.8858, 289.9788, 289.9211, 
    289.9095, 290.0029, 290.1379, 290.1317, 290.0609, 290.1707, 290.1514, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.2688, 287.7101, 
    287.0376, 287.9911, 289.4006, 289.374, 289.1331, 289.2959, 289.4165, 
    289.7666, 289.779, 289.8736, 290.092, 290.1815, 290.0183, 290.1343, 
    289.0108, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.0235, 287.7717, 
    288.2054, 288.9861, 289.1641, 288.7451, 288.5554, 289.0693, 289.5652, 
    289.6047, 289.6833, 289.7623, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 289.0414, _, _, 
    289.0278, 288.9343, 288.8988, 288.5019, 288.4725, 289.0719, 289.4144, 
    289.3297, 289.256, 289.3869, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.4372, 
    288.2567, 288.0349, 288.3616, 289.0509, 289.2039, 289.0234, 288.9597, 
    286.6048, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.2201, 
    287.6134, 287.6531, 287.7771, 288.8992, 289.0154, 288.6852, 288.6726, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 288.9832, 
    287.3656, 287.091, 287.6107, 288.597, 288.5992, 288.4672, 288.4631, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 286.5033, 286.5078, 286.5589, 286.4059, 
    286.2843, 286.8953, _, _, 287.1081, _, _, 287.0089, 287.0491, 286.9807, 
    286.8501, 287.9355, 288.326, 288.1209, 288.283, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 286.2656, 286.3954, 286.0769, 286.5435, 286.6902, 
    286.4923, 286.8853, _, _, _, _, _, 287.0887, 286.7137, 286.6192, 
    286.6214, 288.1745, 288.889, 288.4898, 288.4035, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 285.9996, 285.8991, 285.7099, 286.1579, 286.4685, 
    286.4188, 286.6927, _, _, _, _, _, 287.399, 287.0774, 286.6483, 286.7783, 
    288.305, 289.0052, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 286.1573, 286.0478, 286.2798, 286.3049, 
    286.5372, 290.865, _, 286.1756, 285.7912, 286.1209, 286.8052, 287.1951, 
    287.1326, 286.9729, 287.469, 288.3956, 288.7322, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, 286.4374, 286.8059, 286.1105, 286.663, _, _, 
    286.3257, 285.7816, 286.0656, 286.34, 286.2941, 286.6494, 286.8855, 
    287.3857, 288.0539, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.4637, _, _, 286.1945, 
    286.0993, 286.183, 285.9071, 286.584, 286.88, 287.0893, 287.8431, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.4201, 286.3463, 286.4342, 
    286.3056, 286.2838, 286.5543, 286.6698, 286.7039, 286.9852, 287.4958, 
    287.8153, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 286.1508, _, 285.9833, 285.9005, 
    286.0808, 286.2644, 286.6368, 286.9926, 287.0126, 287.2204, 282.9828, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.4563, 284.8804, 285.4313, 
    285.7052, 286.2932, 286.7198, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.534, 285.5797, 285.1453, 
    283.9334, 284.2205, 284.976, 285.6287, 285.9734, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 286.7185, 286.348, 285.5017, 
    284.6008, 283.6218, 283.6934, 284.1864, 285.1573, 285.8832, 286.7829, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.8824, 285.3122, 284.0973, 
    283.4314, 283.4071, 283.5967, 284.2269, 284.7145, 285.1523, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.9226, 283.6091, 284.4514, 
    284.2624, 283.8799, 283.4893, 284.1117, 285.1955, 286.0553, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 286.7564, 285.0355, 284.1194, 
    284.1986, 284.7971, 284.936, 285.0464, 285.113, 285.5502, 286.2866, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 288.301, _, 286.5396, 285.2831, 285.2737, 
    284.602, 284.2742, 285.082, 285.8584, 286.2307, 286.3463, 286.2835, 
    286.5227, 285.5582, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 285.3004, _, 285.2621, _, 286.619, 
    285.0659, 284.5543, 284.7871, 286.0163, 287.0072, 285.2676, 287.2591, 
    286.8535, 285.9545, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 286.7868, 285.2153, _, _, 285.0043, 
    285.6335, 284.7318, 284.6591, 285.3801, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 285.4144, 287.6729, _, _, 284.999, 
    285.3437, 284.9698, 285.2315, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 285.4602, 285.3091, _, _, 285.4135, 
    285.3999, 285.312, 285.3773, 285.2191, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.0319, 285.2554, 
    285.8444, 285.8252, 289.3625, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.4642, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.149, 
    286.7287, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    285.0882, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    284.1476, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    283.7658, 283.1052, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 287.0961, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 282.4529, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.3916, 285.7069, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.9626, 285.4392, 285.1649, 
    284.8599, 285.3223, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.44, 284.9334, 284.4516, 
    284.6942, 284.3931, 284.677, 284.355, 284.6339, 284.4707, 284.3437, 
    283.656, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.4002, 284.6782, 
    284.2795, 284.3771, 284.4537, 284.4914, 284.4737, 284.5879, 284.619, 
    284.2422, 284.1758, 284.0728, 284.0857, 284.265, 281.9311, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.9406, 284.7485, 
    284.5226, 284.3928, 284.342, 284.2387, 284.2326, 284.3346, 284.1154, 
    284.0941, 283.9278, 284.1088, 284.2519, 284.5482, 285.0346, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.5917, 
    284.0804, 284.1877, 284.0894, 283.9026, 283.9589, 283.8931, 283.9208, 
    283.8269, 283.9123, 284.2851, 284.6748, 285.281, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 285.6174, 283.2317, 
    283.338, 283.7887, 283.8638, 283.7563, 283.7133, 283.7673, 283.7096, 
    283.6598, 283.7292, 283.8495, 284.2229, 284.7439, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.629, 284.9067, 284.3394, 
    283.5785, 283.0178, 283.2771, 283.3976, 283.4997, 283.4326, 283.3812, 
    283.4995, 283.5133, 283.4118, 283.4095, 283.5427, 283.8365, 284.4814, 
    282.5584, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.3105, 284.9644, 284.1908, 
    283.6443, 282.8962, 282.8759, 283.1303, 283.0677, 283.3294, 283.1593, 
    283.2867, 283.2705, 283.2184, 283.1651, 283.3048, 283.4277, 283.7771, 
    284.5127, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.7072, 282.8708, 
    282.6124, 282.8806, 282.9864, 283.2241, 283.1862, 283.1607, 283.0788, 
    283.0941, 283.0787, 283.1272, 283.1694, 283.1752, 283.7955, 284.493, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.4801, 282.774, 
    282.621, 282.7203, 282.8988, 283.086, 283.1407, 283.1137, 283.0104, 
    282.9919, 282.9883, 282.9923, 283.0225, 283.1411, 283.6007, 284.2275, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.4458, 282.4614, 
    282.618, 283.0696, 282.9595, 282.9907, 283.0844, 283.0688, 283.0089, 
    282.9771, 282.9734, 283.0378, 283.148, 283.2076, 283.5492, 284.2852, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.9515, 283.3659, 
    282.3213, 282.5727, 283.0559, 282.9279, 282.8856, 282.8787, 282.8456, 
    282.9978, 283.0226, 283.0483, 283.2609, 283.3362, 283.5026, 284.0437, 
    283.4649, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.6381, 283.0281, 
    282.9072, 283.0018, 283.0231, 282.8636, 282.5173, 282.687, 282.9584, 
    283.0473, 283.1559, 283.4531, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 284.7537, _, _, 
    283.5863, 283.1584, 283.0362, 282.7862, 282.5762, 282.7491, 282.9301, 
    283.019, 283.2259, 283.4978, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.7362, 
    282.5888, 282.453, 282.4656, 282.7751, 282.8607, 282.9716, 283.3833, 
    282.1847, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.9133, 
    282.4411, 282.1886, 282.2112, 282.7979, 282.8334, 282.9146, 283.4636, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.3785, 
    282.37, 281.8863, 282.2094, 282.7378, 282.7118, 282.9731, 283.399, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 283.0818, 283.0296, 283.0663, 282.9987, 
    283.0744, 283.9388, _, _, 283.7025, _, _, 282.5488, 282.2417, 281.8681, 
    281.739, 282.4269, 282.5919, 282.5378, 283.0493, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 282.9465, 283.0042, 282.6276, 282.9671, 283.1214, 
    283.1075, 283.7814, _, _, _, _, _, 282.5915, 281.945, 281.4537, 281.5175, 
    282.4682, 282.9406, 282.9764, 283.3282, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 282.6429, 282.5435, 282.386, 282.6242, 282.8622, 
    283.0226, 283.4593, _, _, _, _, _, 282.7028, 282.1367, 281.4933, 
    281.6445, 282.5317, 283.1124, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 282.7012, 282.638, 282.7393, 282.7311, 283.1116, 
    284.4904, _, 281.9365, 281.7416, 281.8726, 282.2731, 282.4114, 282.0591, 
    281.6619, 281.9588, 282.6848, 283.0117, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, 283.0309, 283.2704, 282.6825, 283.3315, _, _, 
    282.0031, 281.7551, 281.6701, 281.6452, 281.4671, 281.5367, 281.4598, 
    281.8354, 282.5799, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.4009, _, _, 282.0402, 
    281.5789, 281.5163, 281.1196, 281.3399, 281.3721, 281.7532, 282.6159, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.3323, 282.3973, 282.2494, 
    281.8924, 281.5558, 281.6249, 281.5374, 281.3497, 281.5652, 282.2935, 
    282.882, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 283.0839, _, 281.9324, 281.5443, 
    281.423, 281.3465, 281.4381, 281.5503, 281.6444, 282.093, 280.6955, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.3969, 280.9151, 281.0381, 
    280.9125, 281.1339, 281.4516, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.6441, 281.8491, 281.0755, 
    279.9936, 279.781, 280.2499, 280.7155, 281.13, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 283.395, 281.6608, 281.9125, 
    280.8885, 279.8352, 279.4917, 279.6544, 280.2109, 280.7488, 282.2155, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.0133, 281.8979, 280.7276, 
    279.8468, 279.4764, 279.3244, 279.6036, 279.7881, 280.376, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.282, 280.4339, 280.6869, 
    280.3646, 279.7093, 279.2992, 279.6254, 280.3089, 281.2672, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.3654, 281.8959, 280.9109, 
    280.6649, 280.8914, 280.8453, 280.7086, 280.5747, 280.7263, 281.4169, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 283.3604, _, 281.8822, 282.334, 282.0959, 
    281.3579, 280.9196, 281.2815, 281.7544, 281.9246, 281.8266, 281.6235, 
    281.712, 283.4865, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 282.2896, _, 282.7019, _, 281.9774, 
    281.9068, 281.0817, 281.0488, 281.9063, 282.6428, 282.9193, 282.7767, 
    282.1606, 281.2916, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 282.3387, 282.8446, _, _, 282.4884, 
    282.4259, 281.3308, 280.9018, 281.7471, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 281.374, 282.7673, _, _, 282.528, 
    281.9554, 281.2161, 281.2023, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 281.4191, 282.7834, _, _, 282.8824, 
    282.038, 281.724, 281.5378, 281.339, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.1147, 281.4703, 
    282.1198, 282.0717, 284.2584, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 281.9023, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.0648, 
    282.3474, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    281.9962, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    281.3982, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    281.1309, 280.7136, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 282.6024, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 275.9784, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.0114, 279.3362, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 280.3956, 278.9044, 278.3585, 
    278.4568, 279.4353, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.3541, 278.8083, 
    278.4998, 278.9209, 280.776, 278.481, 278.2204, 278.4064, 279.1336, 
    278.7485, 277.7398, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.2802, 278.6844, 
    278.5758, 278.8058, 278.7305, 278.6105, 278.5771, 278.6791, 278.9692, 
    278.8342, 278.7558, 278.6812, 278.776, 278.9861, 275.6859, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.2155, 279.1951, 
    278.9522, 278.6418, 278.6198, 278.7131, 278.7559, 278.8689, 278.8826, 
    279.0459, 279.0084, 279.1171, 279.2147, 279.4004, 280.218, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.6626, 
    278.4621, 278.6301, 278.6469, 278.5466, 278.6327, 278.6881, 278.8656, 
    278.9429, 279.1701, 279.4793, 279.8581, 280.5824, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.349, 277.4847, 
    277.8305, 278.3161, 278.5143, 278.5233, 278.534, 278.6385, 278.6797, 
    278.7825, 278.9913, 279.1873, 279.5336, 280.0423, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.6934, 278.7769, 277.798, 
    277.6465, 277.4601, 277.9289, 278.221, 278.3732, 278.3788, 278.3815, 
    278.5885, 278.7122, 278.7712, 278.8835, 279.057, 279.3043, 279.8828, 
    276.5265, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.6508, 279.1485, 278.2439, 
    277.7754, 277.2811, 277.5834, 278.0277, 278.1198, 278.3702, 278.2985, 
    278.5535, 278.6835, 278.7968, 278.8599, 279.0128, 279.1293, 279.3673, 
    280.0872, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.9056, 277.2305, 
    277.3809, 277.8615, 278.1093, 278.3379, 278.3949, 278.5213, 278.6229, 
    278.8259, 278.9378, 279.0357, 279.1021, 279.195, 279.6837, 280.4549, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.5289, 277.1654, 
    277.3083, 277.7085, 278.0725, 278.2649, 278.3914, 278.5221, 278.6332, 
    278.8463, 279.0091, 279.0708, 279.1293, 279.254, 279.6157, 280.2817, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.3536, 276.9241, 
    277.426, 278.1396, 278.1772, 278.1753, 278.3254, 278.4863, 278.6892, 
    278.9134, 279.0799, 279.2608, 279.4232, 279.4854, 279.7756, 280.5436, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 278.0912, 277.2716, 
    276.6799, 277.3058, 278.0384, 278.0948, 277.9754, 278.1014, 278.2399, 
    278.6755, 278.9628, 279.1833, 279.6146, 279.7414, 279.9819, 280.5683, 
    279.5112, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.554, 277.2837, 
    277.5508, 277.9146, 278.0111, 277.858, 277.841, 278.1685, 278.6107, 
    278.9195, 279.1962, 279.7484, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 279.3675, _, _, 
    278.3523, 278.1007, 277.9303, 277.7931, 277.8475, 278.2489, 278.6031, 
    278.8385, 279.2433, 279.7502, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.699, 
    277.8436, 277.6272, 277.8286, 278.2999, 278.5455, 278.7555, 279.3581, 
    277.3876, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.8669, 
    277.5849, 277.3859, 277.5403, 278.2502, 278.4658, 278.6364, 279.3839, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.7981, 
    277.2483, 277.0132, 277.3859, 278.0191, 278.2356, 278.6688, 279.2542, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 276.6284, 276.5436, 276.5605, 276.5141, 
    276.7373, 278.1476, _, _, 278.8134, _, _, 276.4025, 276.8726, 276.8791, 
    276.7324, 277.3434, 277.7072, 277.9482, 278.7798, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, 276.6301, 276.584, 276.2941, 276.52, 276.6376, 
    276.7683, 277.9614, _, _, _, _, _, 276.9265, 276.7381, 276.433, 276.4041, 
    277.368, 278.0575, 278.4953, 279.1874, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, 276.4303, 276.2627, 276.1474, 276.3459, 276.6057, 
    276.9525, 277.631, _, _, _, _, _, 276.9818, 276.7988, 276.3277, 276.3525, 
    277.3532, 278.3307, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, 276.4069, 276.3329, 276.5137, 276.7322, 
    277.3456, 279.209, _, 275.6004, 275.9927, 276.3754, 276.5535, 276.9289, 
    276.8199, 276.5151, 276.7296, 277.629, 278.2226, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, 277.0319, 277.4233, 277.1527, 278.1513, _, _, 
    276.1138, 276.1121, 276.2096, 276.3955, 276.4879, 276.5175, 276.4657, 
    276.7634, 277.7325, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.2407, _, _, 276.1526, 
    275.9579, 275.972, 275.7936, 276.2259, 276.4047, 276.8011, 277.8921, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.4399, 276.2592, 276.1696, 
    276.0901, 275.961, 276.0767, 276.1452, 276.2087, 276.5672, 277.3601, 
    278.2393, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 277.9302, _, 276.1193, 275.9442, 
    275.8741, 275.9049, 276.0987, 276.3365, 276.6142, 277.1945, 276.2273, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.0761, 275.3687, 275.472, 
    275.5056, 275.9417, 276.6078, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.835, 275.123, 274.774, 
    274.3813, 274.1144, 274.8127, 275.3678, 275.8413, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 277.7208, 276.5618, 275.317, 
    274.3812, 273.5011, 273.4434, 273.9676, 274.7885, 275.4447, 276.211, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.8279, 275.2171, 273.8244, 
    273.0017, 273.0576, 273.2565, 273.9604, 274.6133, 275.0829, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.131, 273.239, 273.5733, 
    273.6579, 273.2554, 272.826, 273.5183, 274.6504, 275.8818, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.4449, 274.8611, 273.8333, 
    273.5907, 273.8875, 273.9905, 273.9485, 274.0675, 274.7556, 275.8722, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 277.2476, _, 276.8729, 275.8372, 275.1948, 
    274.2753, 273.7931, 274.1237, 274.6359, 275.061, 275.2017, 275.5214, 
    276.1702, 278.7335, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 275.8135, _, 276.8533, _, 276.9386, 
    274.9361, 274.0444, 274.175, 275.0705, 275.9094, 277.196, 276.5701, 
    276.7868, 276.184, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 277.6106, 277.1425, _, _, 276.9539, 
    275.53, 274.5593, 274.397, 276.6596, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 275.1494, 277.4685, _, _, 276.7501, 
    275.5091, 274.782, 274.9536, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 275.4593, 277.0785, _, _, 277.411, 
    275.6238, 275.4022, 275.4424, 275.5503, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.9155, 276.117, 
    276.1922, 276.5184, 278.2589, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 276.8246, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 277.5382, 
    277.7264, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    277.5712, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.4272, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    276.3208, 275.9348, _, _, _, _, _, _, _, _, _, _, _, _ ;

 transverse_mercator = _ ;

 time_bnds =
  -173520, -172800,
  -172800, -172080,
  -172080, -171360,
  -171360, -170640,
  -170640, -169920,
  -169920, -169200,
  -169200, -168480,
  -168480, -167760,
  -167760, -167040,
  -167040, -166320,
  -166320, -165600,
  -165600, -164880 ;

 latitude =
  48.8334819352858, 48.8565855874601, 48.8787072756788, 48.899844033934, 
    48.9199930221292, 48.9391515272862, 48.9573169647026, 48.9744868790598, 
    48.9906589454791, 49.005830970526, 49.0200008931604, 49.0331667856326, 
    49.0453268543238, 49.0564794405303, 49.0666230211903, 49.0757562095532, 
    49.0838777557897, 49.0909865475435, 49.0970816104219, 49.1021621084277, 
    49.1062273443289, 49.1092767599682, 49.1113099365105, 49.1123265946288, 
    49.1123265946288, 49.1113099365105, 49.1092767599682, 49.1062273443289, 
    49.1021621084277, 49.0970816104219, 49.0909865475435, 49.0838777557897, 
    49.0757562095532, 49.0666230211903, 49.0564794405303, 49.0453268543238, 
    49.0331667856326, 49.0200008931604, 49.005830970526,
  49.0561868396365, 49.0794714103118, 49.1017664852813, 49.1230690549535, 
    49.1433762374097, 49.1626852796396, 49.1809935587278, 49.1982985829881, 
    49.2145979930463, 49.2298895628688, 49.2441712007369, 49.2574409501642, 
    49.2696969907589, 49.2809376390268, 49.2911613491168, 49.3003667135066, 
    49.3085524636285, 49.3157174704341, 49.3218607448985, 49.3269814384621, 
    49.3310788434097, 49.3341523931884, 49.3362016626606, 49.3372263682953, 
    49.3372263682953, 49.3362016626606, 49.3341523931884, 49.3310788434097, 
    49.3269814384621, 49.3218607448985, 49.3157174704341, 49.3085524636285, 
    49.3003667135066, 49.2911613491168, 49.2809376390268, 49.2696969907589, 
    49.2574409501642, 49.2441712007369, 49.2298895628688,
  49.2788632833994, 49.3023303728217, 49.3248003719413, 49.3462702267173, 
    49.366737012575, 49.3861979356718, 49.4046503341129, 49.4220916791139, 
    49.4385195761098, 49.45393176581, 49.4683261251956, 49.4817006684614, 
    49.4940535478982, 49.5053830547168, 49.5156876198123, 49.5249658144666, 
    49.5332163509902, 49.5404380833014, 49.546630007443, 49.5517912620352, 
    49.5559211286649, 49.5590190322108, 49.5610845411035, 49.5621173675216, 
    49.5621173675216, 49.5610845411035, 49.5590190322108, 49.5559211286649, 
    49.5517912620352, 49.546630007443, 49.5404380833014, 49.5332163509902, 
    49.5249658144666, 49.5156876198123, 49.5053830547168, 49.4940535478982, 
    49.4817006684614, 49.4683261251956, 49.45393176581,
  49.5015109420686, 49.5251621773549, 49.5478086639084, 49.5694473023495, 
    49.5900751245913, 49.6096892951374, 49.6282871123271, 49.6458660095268, 
    49.6624235562675, 49.6779574593248, 49.6924655637426, 49.7059458537976, 
    49.7183964539048, 49.7298156294617, 49.740201787632, 49.7495534780661, 
    49.7578693935594, 49.7651483706457, 49.7713893901275, 49.7765915775401, 
    49.7807542035512, 49.7838766842941, 49.7859585816347, 49.7869996033719, 
    49.7869996033719, 49.7859585816347, 49.7838766842941, 49.7807542035512, 
    49.7765915775401, 49.7713893901275, 49.7651483706457, 49.7578693935594, 
    49.7495534780661, 49.740201787632, 49.7298156294617, 49.7183964539048, 
    49.7059458537976, 49.6924655637426, 49.6779574593248,
  49.724129484382, 49.7479665200925, 49.7707910838008, 49.7926000298754, 
    49.8133903458387, 49.8331591536966, 49.8519037112144, 49.869621413139, 
    49.8863097923637, 49.9019665210362, 49.9165894116077, 49.9301764178223, 
    49.9427256356446, 49.9542353041266, 49.96470380621, 49.9741296694663, 
    49.9825115667709, 49.9898483169126, 49.996138885137, 50.0013823836224, 
    50.0055780718903, 50.0087253571464, 50.0108237945548, 50.0118730874441, 
    50.0118730874441, 50.0108237945548, 50.0087253571464, 50.0055780718903, 
    50.0013823836224, 49.996138885137, 49.9898483169126, 49.9825115667709, 
    49.9741296694663, 49.96470380621, 49.9542353041266, 49.9427256356446, 
    49.9301764178223, 49.9165894116077, 49.9019665210362,
  49.94671857212, 49.9707430908448, 49.9937473484332, 50.0157281520646, 
    50.0366824439681, 50.056607302785, 50.0754999448775, 50.0933577255805, 
    50.1101781403968, 50.1259588261327, 50.1406975619738, 50.1543922704994, 
    50.1670410186342, 50.1786420185368, 50.1891936284237, 50.1986943533267, 
    50.2071428457862, 50.2145379064749, 50.220878484756, 50.2261636791716, 
    50.230392737863, 50.2335650589214, 50.2356801906687, 50.236737831869, 
    50.236737831869, 50.2356801906687, 50.2335650589214, 50.230392737863, 
    50.2261636791716, 50.220878484756, 50.2145379064749, 50.2071428457862, 
    50.1986943533267, 50.1891936284237, 50.1786420185368, 50.1670410186342, 
    50.1543922704994, 50.1406975619738, 50.1259588261327,
  50.1692778598971, 50.1934915728591, 50.2166771686405, 50.238831406269, 
    50.2599511817533, 50.2800335294803, 50.2990756235563, 50.3170747790913, 
    50.3340284534235, 50.3499342472846, 50.364789905903, 50.378593320044, 
    50.3913425269861, 50.4030357114325, 50.4136712063557, 50.4232474937758, 
    50.4317632054701, 50.4392171236146, 50.4456081813557, 50.4509354633116, 
    50.4551982060035, 50.4583957982155, 50.460527781283, 50.4615938493091, 
    50.4615938493091, 50.460527781283, 50.4583957982155, 50.4551982060035, 
    50.4509354633116, 50.4456081813557, 50.4392171236146, 50.4317632054701, 
    50.4232474937758, 50.4136712063557, 50.4030357114325, 50.3913425269861, 
    50.378593320044, 50.364789905903, 50.3499342472846,
  50.3918069949467, 50.4162116426205, 50.4395802490942, 50.4619095242549, 
    50.4831963169386, 50.5034376163633, 50.5226305535041, 50.5407724024097, 
    50.557860581459, 50.5738926545558, 50.5888663322603, 50.6027794728565, 
    50.6156300833537, 50.6274163204212, 50.6381364912556, 50.6477890543787, 
    50.6563726203658, 50.6638859525043, 50.6703279673799, 50.6756977353913, 
    50.6799944811929, 50.683217584064, 50.6853665782046, 50.6864411529576, 
    50.6864411529576, 50.6853665782046, 50.683217584064, 50.6799944811929, 
    50.6756977353913, 50.6703279673799, 50.6638859525043, 50.6563726203658, 
    50.6477890543787, 50.6381364912556, 50.6274163204212, 50.6156300833537, 
    50.6027794728565, 50.5888663322603, 50.5738926545558,
  50.6143056168986, 50.6389029696468, 50.6624562881138, 50.6849622320299, 
    50.7064176020806, 50.7268193413753, 50.7461645368579, 50.7644504206572, 
    50.7816743713754, 50.7978339153141, 50.8129267276349, 50.8269506334545, 
    50.8399036088724, 50.8517837819297, 50.8625894334995, 50.8723189981055, 
    50.8809710646697, 50.8885443771877, 50.895037835331, 50.900450494975, 
    50.9047815686534, 50.9080304259372, 50.9101965937382, 50.9112797565374, 
    50.9112797565374, 50.9101965937382, 50.9080304259372, 50.9047815686534, 
    50.900450494975, 50.895037835331, 50.8885443771877, 50.8809710646697, 
    50.8723189981055, 50.8625894334995, 50.8517837819297, 50.8399036088724, 
    50.8269506334545, 50.8129267276349, 50.7978339153141,
  50.8367733575493, 50.8615652162758, 50.8853049774706, 50.9079892496637, 
    50.9296147843849, 50.9501784776694, 50.9696773715054, 50.9881086552186, 
    51.005469666795, 51.0217578941378, 51.0369709762592, 51.051106704403, 
    51.0641630231004, 51.0761380311534, 51.0870299825486, 51.0968372872976, 
    51.1055585122046, 51.1131923815593, 51.1197377777551, 51.1251937418318, 
    51.1295594739412, 51.1328343337368, 51.135017840685, 51.1361096743002, 
    51.1361096743002, 51.135017840685, 51.1328343337368, 51.1295594739412, 
    51.1251937418318, 51.1197377777551, 51.1131923815593, 51.1055585122046, 
    51.0968372872976, 51.0870299825486, 51.0761380311534, 51.0641630231004, 
    51.051106704403, 51.0369709762592, 51.0217578941378,
  51.0592098406245, 51.0841980374459, 51.1081260021863, 51.1309902911033, 
    51.1527876055376, 51.1735147934582, 51.1931688509468, 51.2117469236191, 
    51.2292463079809, 51.2456644527191, 51.2609989599237, 51.2752475862411, 
    51.2884082439565, 51.3004790020045, 51.3114580869063, 51.3213438836329, 
    51.3301349363928, 51.3378299493437, 51.3444277872271, 51.3499274759254, 
    51.3543282029401, 51.3576293177918, 51.3598303323402, 51.3609309210246, 
    51.3609309210246, 51.3598303323402, 51.3576293177918, 51.3543282029401, 
    51.3499274759254, 51.3444277872271, 51.3378299493437, 51.3301349363928, 
    51.3213438836329, 51.3114580869063, 51.3004790020045, 51.2884082439565, 
    51.2752475862411, 51.2609989599237, 51.2456644527191,
  51.2816146815332, 51.3068010804687, 51.3309190403237, 51.3539650639809, 
    51.3759358015304, 51.396828051855, 51.4166387641529, 51.4353650393964, 
    51.4530041317238, 51.469553449764, 51.4850105578908, 51.4993731774072, 
    51.5126391876562, 51.5248066270584, 51.5358736940742, 51.5458387480901, 
    51.5547003102277, 51.5624570640743, 51.5691078563346, 51.5746516974029, 
    51.5790877618541, 51.5824153888545, 51.5846340824906, 51.5857435120158, 
    51.5857435120158, 51.5846340824906, 51.5824153888545, 51.5790877618541, 
    51.5746516974029, 51.5691078563346, 51.5624570640743, 51.5547003102277, 
    51.5458387480901, 51.5358736940742, 51.5248066270584, 51.5126391876562, 
    51.4993731774072, 51.4850105578908, 51.469553449764,
  51.503987487114, 51.5293739847947, 51.5536837627704, 51.5769132694162, 
    51.5990591024803, 51.6201180107103, 51.6400868954166, 51.6589628119687, 
    51.6767429712244, 51.693424740889, 51.7090056468038, 51.723483374161, 
    51.736855768645, 51.7491208374975, 51.7602767505053, 51.7703218409114, 
    51.7792546062445, 51.7870737090707, 51.7937779776618, 51.7993664065838, 
    51.8038381572005, 51.8071925580963, 51.8094291054129, 51.8105474631041, 
    51.8105474631041, 51.8094291054129, 51.8071925580963, 51.8038381572005, 
    51.7993664065838, 51.7937779776618, 51.7870737090707, 51.7792546062445, 
    51.7703218409114, 51.7602767505053, 51.7491208374975, 51.736855768645, 
    51.723483374161, 51.7090056468038, 51.693424740889,
  51.726327855372, 51.7519163817698, 51.7764198330154, 51.7998346018116, 
    51.8221572324424, 51.8433844224425, 51.8635130242009, 51.882540046498, 
    51.9004626559718, 51.9172781785144, 51.932984100594, 51.9475780705031, 
    51.9610578995302, 51.9734215630539, 51.9846672015575, 51.9947931215643, 
    52.0037977964903, 52.0116798674159, 52.0184381437728, 52.0240716039481, 
    52.0285793958023, 52.0319608371029, 52.0342154158712, 52.0353427906432, 
    52.0353427906432, 52.0342154158712, 52.0319608371029, 52.0285793958023, 
    52.0240716039481, 52.0184381437728, 52.0116798674159, 52.0037977964903, 
    51.9947931215643, 51.9846672015575, 51.9734215630539, 51.9610578995302, 
    51.9475780705031, 51.932984100594, 51.9172781785144,
  51.9486353752078, 51.9744278943847, 51.9991269069176, 52.0227287486397, 
    52.045229909217, 52.0666270338621, 52.0869169249805, 52.1060965437484, 
    52.1241630116184, 52.1411136117533, 52.156945790384, 52.1716571580913, 
    52.1852454910095, 52.1977087319499, 52.2090449914435, 52.2192525487017, 
    52.2283298524923, 52.2362755219323, 52.2430883471937, 52.2487672901243, 
    52.2533114847801, 52.2567202378703, 52.2589930291144, 52.2601295115094, 
    52.2601295115094, 52.2589930291144, 52.2567202378703, 52.2533114847801, 
    52.2487672901243, 52.2430883471937, 52.2362755219323, 52.2283298524923, 
    52.2192525487017, 52.2090449914435, 52.1977087319499, 52.1852454910095, 
    52.1716571580913, 52.156945790384, 52.1411136117533,
  52.1709096261356, 52.1969081370144, 52.2218046324666, 52.2455953902244, 
    52.2682768441492, 52.2898455859909, 52.3102983670786, 52.3296320999401, 
    52.3478438598492, 52.364930886297, 52.3808905843876, 52.3957205261547, 
    52.4094184517975, 52.4219822708356, 52.4334100631803, 52.4437000801209, 
    52.4528507452259, 52.460860655157, 52.467728580395, 52.4734534658772, 
    52.4780344315446, 52.4814707728, 52.4837619608739, 52.4849076431004, 
    52.4849076431004, 52.4837619608739, 52.4814707728, 52.4780344315446, 
    52.4734534658772, 52.467728580395, 52.460860655157, 52.4528507452259, 
    52.4437000801209, 52.4334100631803, 52.4219822708356, 52.4094184517975, 
    52.3957205261547, 52.3808905843876, 52.364930886297,
  52.3931501779927, 52.4193567151496, 52.444452649535, 52.4684341995137, 
    52.4912977419219, 52.5130398138736, 52.533657114497, 52.5531465065976, 
    52.5715050182473, 52.5887298442962, 52.6048183478063, 52.6197680614038, 
    52.6335766885497, 52.6462421047258, 52.6577623585362, 52.6681356727206, 
    52.6773604450806, 52.6854352493164, 52.6923588357728, 52.6981301320942, 
    52.7027482437878, 52.7062124546937, 52.7085222273613, 52.7096772033332, 
    52.7096772033332, 52.7085222273613, 52.7062124546937, 52.7027482437878, 
    52.6981301320942, 52.6923588357728, 52.6854352493164, 52.6773604450806, 
    52.6681356727206, 52.6577623585362, 52.6462421047258, 52.6335766885497, 
    52.6197680614038, 52.6048183478063, 52.5887298442962,
  52.6153565906382, 52.6417732251177, 52.6670705896216, 52.6912448418444, 
    52.7142923003413, 52.7362094463837, 52.7569929257415, 52.7766395503925, 
    52.7951463001544, 52.8125103242383, 52.8287289427218, 52.8437996479383, 
    52.8577201057832, 52.8704881569329, 52.8821018179763, 52.8925592824572, 
    52.9018589218259, 52.9099992862996, 52.9169791056291, 52.9227972897728, 
    52.9274529294748, 52.9309452967488, 52.9332738452656, 52.9344382106436, 
    52.9344382106436, 52.9332738452656, 52.9309452967488, 52.9274529294748, 
    52.9227972897728, 52.9169791056291, 52.9099992862996, 52.9018589218259, 
    52.8925592824572, 52.8821018179763, 52.8704881569329, 52.8577201057832, 
    52.8437996479383, 52.8287289427218, 52.8125103242383,
  52.8375284136417, 52.864157253795, 52.8896580755859, 52.9140269746985, 
    52.9372602101151, 52.9593542060217, 52.9803055536396, 53.000111012981, 
    53.0187675145262, 53.03627216082, 53.052622227985, 53.0678151671508, 
    53.0818486057953, 53.0947203489986, 53.1064283806056, 53.1169708642985, 
    53.1263461445745, 53.1345527476306, 53.1415893821523, 53.147454940006, 
    53.1521484968343, 53.1556693125532, 53.1580168317503, 53.1591906839841, 
    53.1591906839841, 53.1580168317503, 53.1556693125532, 53.1521484968343, 
    53.147454940006, 53.1415893821523, 53.1345527476306, 53.1263461445745, 
    53.1169708642985, 53.1064283806056, 53.0947203489986, 53.0818486057953, 
    53.0678151671508, 53.052622227985, 53.03627216082,
  53.0596651859599, 53.0865083783078, 53.1122147213735, 53.1367802474517, 
    53.1602011546219, 53.1824738087067, 53.2035947451528, 53.2235606708356, 
    53.2423684657828, 53.2600151848149, 53.276498059101, 53.2918144976278, 
    53.3059620885786, 53.3189386006227, 53.3307419841107, 53.3413703721769, 
    53.3508220817457, 53.3590956144406, 53.3661896573958, 53.3721030839683, 
    53.3768349543502, 53.3803845160796, 53.382751204451, 53.3839346428228, 
    53.3839346428228, 53.382751204451, 53.3803845160796, 53.3768349543502, 
    53.3721030839683, 53.3661896573958, 53.3590956144406, 53.3508220817457, 
    53.3413703721769, 53.3307419841107, 53.3189386006227, 53.3059620885786, 
    53.2918144976278, 53.276498059101, 53.2600151848149,
  53.2817664356031, 53.3088261657233, 53.3347401317308, 53.3595043011113, 
    53.3831148096735, 53.40556796356, 53.4268602411813, 53.4469882950702, 
    53.4659489536532, 53.4837392229373, 53.5003562881093, 53.5157975150461, 
    53.5300604517331, 53.5431428295895, 53.5550425646983, 53.5657577589398, 
    53.5752867010263, 53.583627867438, 53.5907799232572, 53.596741722901, 
    53.6015123107512, 53.6050909216801, 53.6074769814724, 53.6086701071415, 
    53.6086701071415, 53.6074769814724, 53.6050909216801, 53.6015123107512, 
    53.596741722901, 53.5907799232572, 53.583627867438, 53.5752867010263, 
    53.5657577589398, 53.5550425646983, 53.5431428295895, 53.5300604517331, 
    53.5157975150461, 53.5003562881093, 53.4837392229373,
  53.5038316792885, 53.5311101727293, 53.55723390191, 53.5821987680465, 
    53.6060008432676, 53.6286363726812, 53.6501017763624, 53.6703936512593, 
    53.6895087730148, 53.7074440977002, 53.7241967634604, 53.7397640920666, 
    53.7541435903751, 53.767332951691, 53.7793300570328, 53.7901329762985, 
    53.7997399693305, 53.808149486878, 53.8153601714553, 53.8213708580963, 
    53.8261805750017, 53.8297885440809, 53.8321941813853, 53.8333970974347, 
    53.8333970974347, 53.8321941813853, 53.8297885440809, 53.8261805750017, 
    53.8213708580963, 53.8153601714553, 53.808149486878, 53.7997399693305, 
    53.7901329762985, 53.7793300570328, 53.767332951691, 53.7541435903751, 
    53.7397640920666, 53.7241967634604, 53.7074440977002,
  53.7258604220818, 53.7533599453023, 53.7796956173633, 53.8048632717073, 
    53.8288589153322, 53.8516787309161, 53.8733190788607, 53.8937764992506, 
    53.9130477137265, 53.9311296272684, 53.9480193298875, 53.9637140982229, 
    53.9782113970432, 53.9915088806482, 54.0036043941706, 54.0144959747761, 
    54.0241818527586, 54.0326604525308, 54.0399303935075, 54.0459904908816, 
    54.050839756291, 54.0544773983756, 54.0569028232237, 54.0581156347076, 
    54.0581156347076, 54.0569028232237, 54.0544773983756, 54.050839756291, 
    54.0459904908816, 54.0399303935075, 54.0326604525308, 54.0241818527586, 
    54.0144959747761, 54.0036043941706, 53.9915088806482, 53.9782113970432, 
    53.9637140982229, 53.9480193298875, 53.9311296272684,
  53.9478521570256, 53.9755750183637, 54.0021248534264, 54.0274974263339, 
    54.05168867746, 54.0746947256158, 54.0965118701513, 54.1171365929701, 
    54.1365655604557, 54.1547956253059, 54.1718238282731, 54.1876473998072, 
    54.2022637616, 54.215670528028, 54.2278655074921, 54.238846703652, 
    54.2486123165538, 54.2571607436492, 54.2644905807054, 54.270600622603, 
    54.2754898640229, 54.2791575000198, 54.2816029264815, 54.2828257404746, 
    54.2828257404746, 54.2816029264815, 54.2791575000198, 54.2754898640229, 
    54.270600622603, 54.2644905807054, 54.2571607436492, 54.2486123165538, 
    54.238846703652, 54.2278655074921, 54.215670528028, 54.2022637616, 
    54.1876473998072, 54.1718238282731, 54.1547956253059,
  54.1698063647541, 54.197754915423, 54.2245211749891, 54.2501008366557, 
    54.2744897726336, 54.2976840363871, 54.3196798647945, 54.3404736802208, 
    54.3600620924993, 54.3784419008183, 54.3956100955118, 54.4115638597505, 
    54.4263005711306, 54.439817803159, 54.4521133266319, 54.4631851109056, 
    54.4730313250573, 54.4816503389343, 54.4890407240904, 54.495201254608, 
    54.5001309078049, 54.5038288648246, 54.5062945111097, 54.5075274367576, 
    54.5075274367576, 54.5062945111097, 54.5038288648246, 54.5001309078049, 
    54.495201254608, 54.4890407240904, 54.4816503389343, 54.4730313250573, 
    54.4631851109056, 54.4521133266319, 54.439817803159, 54.4263005711306, 
    54.4115638597505, 54.3956100955118, 54.3784419008183,
  54.3917225130938, 54.4198991482086, 54.4468841361556, 54.4726730975784, 
    54.4972618349404, 54.5206463348336, 54.5428227702021, 54.5637875024734, 
    54.5835370835974, 54.6020682579881, 54.6193779643662, 54.6354633374993, 
    54.6503217098374, 54.663950613042, 54.6763477794049, 54.6875111431567, 
    54.6974388416621, 54.7061292164999, 54.7135808144277, 54.7197923882281, 
    54.7247628974365, 54.7284915089496, 54.7309775975124, 54.7322207460844, 
    54.7322207460844, 54.7309775975124, 54.7284915089496, 54.7247628974365, 
    54.7197923882281, 54.7135808144277, 54.7061292164999, 54.6974388416621, 
    54.6875111431567, 54.6763477794049, 54.663950613042, 54.6503217098374, 
    54.6354633374993, 54.6193779643662, 54.6020682579881,
  54.6136000566501, 54.6420072162843, 54.6692132798904, 54.6952137938601, 
    54.7200044892762, 54.7435812842874, 54.7659402863956, 54.787077794649, 
    54.8069903017404, 54.8256744960053, 54.843127263319, 54.8593456888872, 
    54.8743270589308, 54.8880688622591, 54.9005687917316, 54.9118247456052, 
    54.9218348287649, 54.9305973538365, 54.9381108421795, 54.9443740247597, 
    54.9493858428978, 54.953145448897, 54.9556522065439, 54.9569056914869, 
    54.9569056914869, 54.9556522065439, 54.953145448897, 54.9493858428978, 
    54.9443740247597, 54.9381108421795, 54.9305973538365, 54.9218348287649, 
    54.9118247456052, 54.9005687917316, 54.8880688622591, 54.8743270589308, 
    54.8593456888872, 54.843127263319, 54.8256744960053,
  54.8354384363769, 54.8640786066519, 54.8915081376524, 54.9177224997749, 
    54.9427173510389, 54.9664885395302, 54.9890321057544, 55.0103442848943, 
    55.0304215089687, 55.0492604088905, 55.0668578164185, 55.0832107660021, 
    55.0983164965153, 55.1121724528775, 55.1247762875587, 55.1361258619669, 
    55.1462192477163, 55.1550547277727, 55.1626307974776, 55.1689461654456, 
    55.1739997543371, 55.1777907015036, 55.1803183595053, 55.1815822964993, 
    55.1815822964993, 55.1803183595053, 55.1777907015036, 55.1739997543371, 
    55.1689461654456, 55.1626307974776, 55.1550547277727, 55.1462192477163, 
    55.1361258619669, 55.1247762875587, 55.1121724528775, 55.0983164965153, 
    55.0832107660021, 55.0668578164185, 55.0492604088905,
  55.0572370791323, 55.0861127933387, 55.1137682290145, 55.1401987787642, 
    55.1654000258095, 55.1893677465041, 55.2120979127551, 55.2335866943471, 
    55.2538304611647, 55.2728257853113, 55.2905694431187, 55.3070584170474, 
    55.3222898974721, 55.3362612843512, 55.3489701887777, 55.3604144344079, 
    55.3705920587683, 55.3795013144363, 55.3871406700942, 55.393508811455, 
    55.3986046420581, 55.4024272839346, 55.4049760781404, 55.4062505851564, 
    55.4062505851564, 55.4049760781404, 55.4024272839346, 55.3986046420581, 
    55.393508811455, 55.3871406700942, 55.3795013144363, 55.3705920587683, 
    55.3604144344079, 55.3489701887777, 55.3362612843512, 55.3222898974721, 
    55.3070584170474, 55.2905694431187, 55.2728257853113,
  55.2789953972162, 55.3081092369699, 55.3359930612691, 55.3626421830744, 
    55.3880521090219, 55.4122185420116, 55.4351373837004, 55.4568047368943, 
    55.4772169078371, 55.4963704083923, 55.514261958113, 55.530888486199, 
    55.5462471333366, 55.5603352534181, 55.5731504151401, 55.5846904034759, 
    55.5949532210214, 55.6039370892128, 55.6116404494124, 55.6180619638627, 
    55.6232005165072, 55.6270552136753, 55.6296253846322, 55.6309105819916, 
    55.6309105819916, 55.6296253846322, 55.6270552136753, 55.6232005165072, 
    55.6180619638627, 55.6116404494124, 55.6039370892128, 55.5949532210214, 
    55.5846904034759, 55.5731504151401, 55.5603352534181, 55.5462471333366, 
    55.530888486199, 55.514261958113, 55.4963704083923,
  55.5007127878905, 55.5300673843242, 55.5581821290187, 55.5850522533813, 
    55.610673185619, 55.6350405534037, 55.6581501864381, 55.6799981189193, 
    55.7005805918965, 55.7198940555174, 55.7379351711615, 55.754700813456, 
    55.7701880721711, 55.784394253993, 55.7973168841697, 55.8089537080294, 
    55.819302692368, 55.8283620267032, 55.8361301243949, 55.8426056236283, 
    55.8477873882598, 55.8516745085238, 55.8542663015992, 55.8555623120351, 
    55.8555623120351, 55.8542663015992, 55.8516745085238, 55.8477873882598, 
    55.8426056236283, 55.8361301243949, 55.8283620267032, 55.819302692368, 
    55.8089537080294, 55.7973168841697, 55.784394253993, 55.7701880721711, 
    55.754700813456, 55.7379351711615, 55.7198940555174,
  55.7223886328819, 55.7519866678729, 55.7803349137503, 55.8074285183992, 
    55.8332628296971, 55.8578333982566, 55.8811359800687, 55.9031665390404, 
    55.9239212494223, 55.943396498124, 55.9615888869117, 55.9784952344855, 
    55.9941125784332, 56.0084381770568, 56.0214695110703, 56.0332042851638, 
    56.0436404294345, 56.0527761006798, 56.0606096835523, 56.0671397915733, 
    56.0723652680058, 56.0762851865827, 56.0788988520912, 56.080205800812, 
    56.080205800812, 56.0788988520912, 56.0762851865827, 56.0723652680058, 
    56.0671397915733, 56.0606096835523, 56.0527761006798, 56.0436404294345, 
    56.0332042851638, 56.0214695110703, 56.0084381770568, 55.9941125784332, 
    55.9784952344855, 55.9615888869117, 55.943396498124,
  55.9440222978651, 55.9738665053015, 56.0024508833942, 56.0297704944765, 
    56.0558206041349, 56.0805966840348, 56.1040944146424, 56.1263096878386, 
    56.1472386094213, 56.1668775014902, 56.1852229047122, 56.2022715804623, 
    56.2180205128378, 56.2324669105415, 56.2456082086313, 56.2574420701342, 
    56.267966387521, 56.2771792840402, 56.2850791149089, 56.2916644683588, 
    56.2969341665357, 56.3008872662513, 56.3035230595856, 56.3048410743402, 
    56.3048410743402, 56.3035230595856, 56.3008872662513, 56.2969341665357, 
    56.2916644683588, 56.2850791149089, 56.2771792840402, 56.267966387521, 
    56.2574420701342, 56.2456082086313, 56.2324669105415, 56.2180205128378, 
    56.2022715804623, 56.1852229047122, 56.1668775014902,
  56.1656131319263, 56.1957062990121, 56.2245294918656, 56.2520776851737, 
    56.2783460602095, 56.3033300077425, 56.3270251308429, 56.349427247575, 
    56.3705323935757, 56.3903368245124, 56.4088370184185, 56.4260296779007, 
    56.4419117322152, 56.4564803392099, 56.4697328871288, 56.4816669962763, 
    56.4922805205387, 56.5015715487596, 56.5095384059689, 56.5161796544613, 
    56.521494094725, 56.5254807662164, 56.5281389479827, 56.5294681591286, 
    56.5294681591286, 56.5281389479827, 56.5254807662164, 56.521494094725, 
    56.5161796544613, 56.5095384059689, 56.5015715487596, 56.4922805205387, 
    56.4816669962763, 56.4697328871288, 56.4564803392099, 56.4419117322152, 
    56.4260296779007, 56.4088370184185, 56.3903368245124,
  56.3871604670056, 56.4175054356075, 56.4465701785876, 56.4743495808264, 
    56.5008387371962, 56.5260329555599, 56.5499277596605, 56.5725188918969, 
    56.5938023159816, 56.6137742194748, 56.6324310161924, 56.6497693484814, 
    56.6657860893624, 56.6804783445315, 56.6938434542224, 56.7058789949228, 
    56.7165827809443, 56.7259528658414, 56.7339875436794, 56.7406853501479, 
    56.7460450635182, 56.7500657054437, 56.7527465416015, 56.7540870821748, 
    56.7540870821748, 56.7527465416015, 56.7500657054437, 56.7460450635182, 
    56.7406853501479, 56.7339875436794, 56.7259528658414, 56.7165827809443, 
    56.7058789949228, 56.6938434542224, 56.6804783445315, 56.6657860893624, 
    56.6497693484814, 56.6324310161924, 56.6137742194748,
  56.6086636173186, 56.6392632853541, 56.6685723679967, 56.6965856580905, 
    56.7232981619533, 56.748705102466, 56.7728019220507, 56.7955842855321, 
    56.8170480828776, 56.8371894318102, 56.8560046802916, 56.87349040887, 
    56.8896434328887, 56.9044608045526, 56.9179398148487, 56.9300779953174, 
    56.9408731196724, 56.9503232052652, 56.9584265143936, 56.9651815554507, 
    56.9705870839134, 56.9746421031687, 56.9773458651756, 56.9786978709633, 
    56.9786978709633, 56.9773458651756, 56.9746421031687, 56.9705870839134, 
    56.9651815554507, 56.9584265143936, 56.9503232052652, 56.9408731196724, 
    56.9300779953174, 56.9179398148487, 56.9044608045526, 56.8896434328887, 
    56.87349040887, 56.8560046802916, 56.8371894318102,
  56.8301218787543, 56.8609792016248, 56.8905354690274, 56.9187853794693, 
    56.9457238484902, 56.9713460118464, 56.9956472285803, 57.0186230839715, 
    57.0402693923616, 57.0605821998495, 57.0795577868526, 57.0971926705288, 
    57.1134836070555, 57.1284275937617, 57.14202187111, 57.1542639245252, 
    57.1651514860652, 57.174682535934, 57.1828553038313, 57.1896682701396, 
    57.1951201669444, 57.1992099788869, 57.2019369438483, 57.2033005534631, 
    57.2033005534631, 57.2019369438483, 57.1992099788869, 57.1951201669444, 
    57.1896682701396, 57.1828553038313, 57.174682535934, 57.1651514860652, 
    57.1542639245252, 57.14202187111, 57.1284275937617, 57.1134836070555, 
    57.0971926705288, 57.0795577868526, 57.0605821998495,
  57.0515345282499, 57.0826525203189, 57.1124588745778, 57.1409481928223, 
    57.1681152975183, 57.1939552350846, 57.2184632790585, 57.2416349331383, 
    57.2634659340969, 57.2839522545632, 57.3030901056635, 57.3208759395213, 
    57.3373064516091, 57.352378582949, 57.3660895221587, 57.3784367073389, 
    57.3894178277987, 57.3990308256174, 57.4072738970385, 57.4141454936951, 
    57.4196443236636, 57.4237693523442, 57.4265198031676, 57.4278951581257, 
    57.4278951581257, 57.4265198031676, 57.4237693523442, 57.4196443236636, 
    57.4141454936951, 57.4072738970385, 57.3990308256174, 57.3894178277987, 
    57.3784367073389, 57.3660895221587, 57.352378582949, 57.3373064516091, 
    57.3208759395213, 57.3030901056635, 57.2839522545632,
  57.272900823141, 57.3042825592593, 57.3343419609531, 57.3630735308539, 
    57.3904719959833, 57.4165323111379, 57.4412496621536, 57.4646194690438, 
    57.4866373890061, 57.5072993192908, 57.5266013999282, 57.544540016308, 
    57.5611118016069, 57.5763136390607, 57.5901426640766, 57.6025962661819, 
    57.6136720908064, 57.6233680408944, 57.6316822783454, 57.638613225279, 
    57.6441595651236, 57.6483202435262, 57.651094469082, 57.6524817138827, 
    57.6524817138827, 57.651094469082, 57.6483202435262, 57.6441595651236, 
    57.638613225279, 57.6316822783454, 57.6233680408944, 57.6136720908064, 
    57.6025962661819, 57.5901426640766, 57.5763136390607, 57.5611118016069, 
    57.544540016308, 57.5266013999282, 57.5072993192908,
  57.494220000485, 57.525868617566, 57.5561840872864, 57.5851608105813, 
    57.6127934165797, 57.6390767660954, 57.6640059549939, 57.6875763174304, 
    57.7097834289522, 57.7306231094597, 57.750091426021, 57.7681846955346, 
    57.7848994872367, 57.8002326250469, 57.8141811897497, 57.8267425210072, 
    57.8379142192, 57.8476941470928, 57.8560804313222, 57.8630714637041, 
    57.8686659023583, 57.872862672648, 57.8756609679347, 57.877060250144, 
    57.877060250144, 57.8756609679347, 57.872862672648, 57.8686659023583, 
    57.8630714637041, 57.8560804313222, 57.8476941470928, 57.8379142192, 
    57.8267425210072, 57.8141811897497, 57.8002326250469, 57.7848994872367, 
    57.7681846955346, 57.750091426021, 57.7306231094597,
  57.7154912763585, 57.7474099750036, 57.7779845949369, 57.8072094327815, 
    57.8350790172446, 57.861588112718, 57.8867317227521, 57.9105050933977, 
    57.9329037164074, 57.9539233322928, 57.9735599332302, 57.9918097658104, 
    58.0086693336277, 58.0241353997031, 58.0382049887377, 58.0508753891916, 
    58.0621441551863, 58.0720091082258, 58.0804683387334, 58.0875202074035, 
    58.0931633463629, 58.097396660143, 58.1002193264589, 58.1016307967947, 
    58.1016307967947, 58.1002193264589, 58.097396660143, 58.0931633463629, 
    58.0875202074035, 58.0804683387334, 58.0720091082258, 58.0621441551863, 
    58.0508753891916, 58.0382049887377, 58.0241353997031, 58.0086693336277, 
    57.9918097658104, 57.9735599332302, 57.9539233322928,
  57.9367138451252, 57.9689058913026, 57.9997428068629, 58.0292187814151, 
    58.057328240631, 58.0840658499596, 58.1094265182131, 58.1334054010153, 
    58.1559979041072, 58.1771996865032, 58.1970066634925, 58.2154150094787, 
    58.2324211606547, 58.2480218175057, 58.2622139471378, 58.2749947854262, 
    58.2863618389813, 58.2963128869272, 58.3048459824905, 58.3119594543972, 
    58.3176519080737, 58.3219222266514, 58.3247695717722, 58.3261933841937, 
    58.3261933841937, 58.3247695717722, 58.3219222266514, 58.3176519080737, 
    58.3119594543972, 58.3048459824905, 58.2963128869272, 58.2863618389813, 
    58.2749947854262, 58.2622139471378, 58.2480218175057, 58.2324211606547, 
    58.2154150094787, 58.1970066634925, 58.1771996865032,
  58.1578868786747, 58.1903556054534, 58.2214580269698, 58.2511882230267, 
    58.2795405135593, 58.3065094624688, 58.3320898813233, 58.3562768329185, 
    58.3790656346907, 58.4004518619769, 58.4204313511149, 58.4390002023768, 
    58.4561547827333, 58.4718917284397, 58.486207947443, 58.4991006216021, 
    58.51056720872, 58.5206054443828, 58.529213343602, 58.536389202259, 
    58.5421315983467, 58.5464393930084, 58.549311731371, 58.5507480431706, 
    58.5507480431706, 58.549311731371, 58.5464393930084, 58.5421315983467, 
    58.536389202259, 58.529213343602, 58.5206054443828, 58.51056720872, 
    58.4991006216021, 58.486207947443, 58.4718917284397, 58.4561547827333, 
    58.4390002023768, 58.4204313511149, 58.4004518619769,
  58.37900952563, 58.4117583349704, 58.4431295394302, 58.4731171061201, 
    58.5017152464466, 58.5289184200693, 58.5547213387214, 58.5791189698868, 
    58.6021065403257, 58.6236795394418, 58.6438337224855, 58.6625651135859, 
    58.6798700086067, 58.69574497782, 58.7101868683945, 58.7231928066908, 
    58.7347602003629, 58.7448867402593, 58.7535704021222, 58.7608094480806, 
    58.766602427935, 58.7709481802318, 58.773845833125, 58.7752948050235, 
    58.7752948050235, 58.773845833125, 58.7709481802318, 58.766602427935, 
    58.7608094480806, 58.7535704021222, 58.7448867402593, 58.7347602003629, 
    58.7231928066908, 58.7101868683945, 58.69574497782, 58.6798700086067, 
    58.6625651135859, 58.6438337224855, 58.6236795394418,
  58.6000809105225, 58.633113275127, 58.664756607977, 58.6950047605081, 
    58.7238518327113, 58.7512921772186, 58.7773204032489, 58.8019313804052, 
    58.8251202423176, 58.8468823901224, 58.8672134957723, 58.8861095051706, 
    58.9035666411234, 58.9195814061045, 58.9341505848275, 58.9472712466204, 
    58.9589407475983, 58.9691567326303, 58.977917137097, 58.985220188435, 
    58.9910644074661, 58.9954486095092, 58.9983719052711, 58.9998337015167, 
    58.9998337015167, 58.9983719052711, 58.9954486095092, 58.9910644074661, 
    58.985220188435, 58.977917137097, 58.9691567326303, 58.9589407475983, 
    58.9472712466204, 58.9341505848275, 58.9195814061045, 58.9035666411234, 
    58.8861095051706, 58.8672134957723, 58.8468823901224,
  58.8211001329322, 58.854419598157, 58.8863384751658, 58.9168504966345, 
    58.9459496481529, 58.9736301724444, 58.9998865734409, 59.0247136202068, 
    59.0481063507023, 59.0700600753805, 59.0905703806082, 59.1096331319069, 
    59.1272444770054, 59.1434008486992, 59.1580989675106, 59.1713358441455, 
    59.1831087817406, 59.193415377899, 59.2022535265081, 59.2096214193382, 
    59.215517547418, 59.2199407021848, 59.2228899764071, 59.2243647648779, 
    59.2243647648779, 59.2228899764071, 59.2199407021848, 59.215517547418, 
    59.2096214193382, 59.2022535265081, 59.193415377899, 59.1831087817406, 
    59.1713358441455, 59.1580989675106, 59.1434008486992, 59.1272444770054, 
    59.1096331319069, 59.0905703806082, 59.0700600753805,
  59.0420662665924, 59.0756764524242, 59.1078743616072, 59.1386536048674, 
    59.168008050306, 59.1959318277561, 59.2224193329944, 59.2474652317953, 
    59.2710644638209, 59.2932122463396, 59.3139040777633, 59.3331357409991, 
    59.3509033066065, 59.3672031357554, 59.3820318829783, 59.3953864987121, 
    59.4072642316239, 59.4176626307174, 59.4265795472143, 59.4340131362092, 
    59.4399618580934, 59.4444244797453, 59.4474000754857, 59.4488880277957, 
    59.4488880277957, 59.4474000754857, 59.4444244797453, 59.4399618580934, 
    59.4340131362092, 59.4265795472143, 59.4176626307174, 59.4072642316239, 
    59.3953864987121, 59.3820318829783, 59.3672031357554, 59.3509033066065, 
    59.3331357409991, 59.3139040777633, 59.2932122463396,
  59.2629783584575, 59.2968829615559, 59.3293634651655, 59.3604133547633, 
    59.3900263777658, 59.4181965480319, 59.4449181502137, 59.4701857439476, 
    59.4939941678764, 59.5163385434936, 59.5372142788027, 59.5566170717837, 
    59.5745429136596, 59.5909880919573, 59.6059491933558, 59.6194231063166, 
    59.6314070234915, 59.6418984439026, 59.6508951748907, 59.6583953338285, 
    59.6643973495945, 59.668899963806, 59.6719022318081, 59.6734035234171, 
    59.6734035234171, 59.6719022318081, 59.668899963806, 59.6643973495945, 
    59.6583953338285, 59.6508951748907, 59.6418984439026, 59.6314070234915, 
    59.6194231063166, 59.6059491933558, 59.5909880919573, 59.5745429136596, 
    59.5566170717837, 59.5372142788027, 59.5163385434936,
  59.4838354277295, 59.5180382235396, 59.5508049601247, 59.582128994298, 
    59.6120039494857, 59.640423720379, 59.667382477432, 59.6928746711945, 
    59.7168950364712, 59.7394385962984, 59.7605006657293, 59.7800768554206, 
    59.7981630750135, 59.814755536301, 59.8298507561769, 59.8434455593584, 
    59.8555370808796, 59.8661227683484, 59.8752003839648, 59.8827680062943, 
    59.8888240317951, 59.8933671760952, 59.8963964750164, 59.8979112853448, 
    59.8979112853448, 59.8963964750164, 59.8933671760952, 59.8888240317951, 
    59.8827680062943, 59.8752003839648, 59.8661227683484, 59.8555370808796, 
    59.8434455593584, 59.8298507561769, 59.814755536301, 59.7981630750135, 
    59.7800768554206, 59.7605006657293, 59.7394385962984,
  59.7046364648451, 59.7391413097821, 59.7721979963169, 59.8037997490664, 
    59.8339400640435, 59.8626127134664, 59.8898117504082, 59.9155315132783, 
    59.9397666301241, 59.9625120227452, 59.9837629106106, 60.0035148145708, 
    60.0217635603576, 60.038505281863, 60.0537364241927, 60.0674537464858, 
    60.079654324497, 60.0903355529345, 60.0994951475502, 60.1071311469774, 
    60.1132419143128, 60.1178261384393, 60.1208828350877, 60.1224113476344, 
    60.1224113476344, 60.1208828350877, 60.1178261384393, 60.1132419143128, 
    60.1071311469774, 60.0994951475502, 60.0903355529345, 60.079654324497, 
    60.0674537464858, 60.0537364241927, 60.038505281863, 60.0217635603576, 
    60.0035148145708, 59.9837629106106, 59.9625120227452,
  59.9253804304179, 59.9601912641265, 59.9935416982147, 60.0254248214456, 
    60.055833998876, 60.0847628768277, 60.1122053876966, 60.1381557545877, 
    60.1626084957663, 60.1855584289152, 60.2070006751896, 60.2269306630599, 
    60.2453441319351, 60.2622371355591, 60.277606045173, 60.2914475524356, 
    60.3037586720989, 60.31453674443, 60.3237794373771, 60.3314847484739, 
    60.3376510064788, 60.3422768727461, 60.3453613423259, 60.3469037447916, 
    60.3469037447916, 60.3453613423259, 60.3422768727461, 60.3376510064788, 
    60.3314847484739, 60.3237794373771, 60.31453674443, 60.3037586720989, 
    60.2914475524356, 60.277606045173, 60.2622371355591, 60.2453441319351, 
    60.2269306630599, 60.2070006751896, 60.1855584289152,
  60.1460662541356, 60.1811871018278, 60.2148351639827, 60.2470033897233, 
    60.2776850094805, 60.3068735401344, 60.3345627899887, 60.360746863566, 
    60.3854201662143, 60.4085774085145, 60.4302136104778, 60.4503241055256, 
    60.468904544242, 60.4859508978922, 60.501459461698, 60.5154268578652, 
    60.5278500383548, 60.5387262873938, 60.54805322372, 60.5558288025559, 
    60.5620513173079, 60.5667194009883, 60.569832027355, 60.5713885117696, 
    60.5713885117696, 60.569832027355, 60.5667194009883, 60.5620513173079, 
    60.5558288025559, 60.54805322372, 60.5387262873938, 60.5278500383548, 
    60.5154268578652, 60.501459461698, 60.4859508978922, 60.468904544242, 
    60.4503241055256, 60.4302136104778, 60.4085774085145 ;

 longitude =
  -10.0099032089996, -9.67231824107548, -9.33431249451303, -8.99590363883535, 
    -8.65710948045695, -8.31794795720088, -7.97843713268945, 
    -7.63859519061489, -7.29844042889601, -6.95799125372699, 
    -6.61726617352461, -6.27628379277987, -5.93506280582035, 
    -5.59362199048939, -5.25198020174822, -4.91015636520727, 
    -4.56816947059276, -4.2260385651548, -3.88378274702307, 
    -3.54142115851636, -3.19897297941198, -2.85645742018132, 
    -2.51389371519774, -2.17130111592281, -1.82869888407719, 
    -1.48610628480226, -1.14354257981868, -0.801027020588025, 
    -0.458578841483637, -0.116217252976927, 0.226038565154795, 
    0.568169470592757, 0.910156365207267, 1.25198020174822, 1.59362199048939, 
    1.93506280582035, 2.27628379277987, 2.61726617352461, 2.95799125372699,
  -10.0458624695909, -9.7067994526941, -9.36730898608934, -9.02740900763868, 
    -8.68711759578541, -8.34645296393427, -8.00543345470023, 
    -7.66407753403265, -7.32240378522081, -6.98043090278747, 
    -6.63817768627677, -6.29566303394286, -5.95290593634568, 
    -5.60992546986037, -5.26674079010657, -4.92337112530408, 
    -4.57983576956137, -4.23615407610318, -3.89234545044372, 
    -3.54842934351185, -3.20442524473469, -2.86035267508588, 
    -2.51623118010518, -2.17208032289559, -1.82791967710441, 
    -1.48376881989482, -1.13964732491413, -0.795574755265315, 
    -0.451570656488147, -0.107654549556285, 0.236154076103178, 
    0.579835769561371, 0.923371125304078, 1.26674079010657, 1.60992546986037, 
    1.95290593634568, 2.29566303394286, 2.63817768627677, 2.98043090278747,
  -10.0822669886824, -9.74170813230963, -9.40071500855603, -9.05930582921149, 
    -8.71749895045653, -8.37531286710161, -8.03276620668996, 
    -7.68987772347056, -7.34666629224811, -7.00315090211636, 
    -6.65935065008181, -6.31528473458406, -5.97097244891979, 
    -5.62643317457679, -5.28168637448489, -4.93675158619024, 
    -4.59164841495978, -4.24639652682248, -3.90101564155395, 
    -3.55552552561118, -3.20994598502401, -2.86429685824996, 
    -2.51859800899918, -2.17286931903601, -1.82713068096399, 
    -1.48140199100082, -1.13570314175004, -0.790054014975992, 
    -0.444474474388818, -0.0989843584460488, 0.246396526822481, 
    0.59164841495978, 0.936751586190235, 1.28168637448489, 1.62643317457679, 
    1.97097244891979, 2.31528473458406, 2.65935065008181, 3.00315090211636,
  -10.1191238541792, -9.77705109793588, -9.43453710606329, -9.0916003700088, 
    -8.74825952954401, -8.40453336685909, -8.06044080051507, 
    -7.7160008792613, -7.37123277572486, -7.02615577997884, 
    -6.68078929299644, -6.33515281999788, -5.98926596369688, 
    -5.64314841745374, -5.296819958342, -4.95030044013536, -4.60360978622214, 
    -4.25676798245379, -3.90979506993475, -3.56271113776034, 
    -3.21553631570961, -2.86829076690028, -2.52099468041237, 
    -2.17366826388774, -1.82633173611226, -1.47900531958763, 
    -1.13170923309972, -0.784463684290387, -0.437288862239664, 
    -0.0902049300652483, 0.256767982453785, 0.603609786222135, 
    0.950300440135361, 1.29681995834199, 1.64314841745374, 1.98926596369687, 
    2.33515281999788, 2.68078929299644, 3.02615577997883,
  -10.1564403101608, -9.81283531816545, -9.46878196761471, -9.1242990354882, 
    -8.77940545115234, -8.4341202903053, -8.0884627687744, -7.74245223617316, 
    -7.39610816942524, -7.04945016616247, -6.70249793800405, 
    -6.35527130372431, -6.00779018231606, -5.66007458595679, 
    -5.31214461288497, -4.96402044019351, -4.61572231654769, 
    -4.26727055483479, -3.91868552475244, -3.56998764534307, 
    -3.22119737748155, -2.87233521632329, -2.52342168371991, 
    -2.17447732060972, -1.82552267939028, -1.4765783162801, 
    -1.12766478367671, -0.778802622518448, -0.430012354656932, 
    -0.0813144752475589, 0.267270554834791, 0.61572231654769, 
    0.964020440193505, 1.31214461288497, 1.66007458595679, 2.00779018231606, 
    2.35527130372431, 2.70249793800405, 3.04945016616247,
  -10.1942237611228, -9.84906791627151, -9.50345643102423, -9.15740837391722, 
    -8.81094297006977, -8.4640795949756, -8.11683776814049, 
    -7.76923714657417, -7.42129751814363, -7.07303879479541, 
    -6.72448100565447, -6.37564429000698, -6.02654889017454, 
    -5.67721514428742, -5.32766347896419, -4.97791440190527, 
    -4.62798849440789, -4.27790640380992, -3.92768883587013, 
    -3.57735654709223, -3.2269303370003, -2.87643104037305, 
    -2.52587951944441, -2.17529665607787, -1.82470334392213, 
    -1.47412048055559, -1.12356895962695, -0.773069662999705, 
    -0.422643452907771, -0.0723111641298666, 0.277906403809922, 
    0.627988494407887, 0.977914401905269, 1.32766347896419, 1.67721514428742, 
    2.02654889017454, 2.37564429000698, 2.72448100565447, 3.07303879479541,
  -10.2324817763575, -9.88575617444401, -9.53856748700325, -9.19093508030624, 
    -8.84287848154239, -8.49441737245244, -8.14557158280176, 
    -7.79636108370186, -7.44680598078773, -7.09692650725897, 
    -6.74674301679238, -6.39627597633386, -6.04554595877738, 
    -5.69457363553879, -5.34337976903234, -4.99198520505758, 
    -4.64041086510456, -4.28867773858492, -3.93680687499694, 
    -3.58481937603209, -3.23273638763094, -2.88057909199631, 
    -2.52836869957134, -2.17612644099025, -1.82387355900975, 
    -1.47163130042867, -1.11942090800369, -0.767263612369062, 
    -0.415180623967913, -0.06319312500306, 0.288677738584914, 
    0.640410865104554, 0.991985205057582, 1.34337976903233, 1.69457363553878, 
    2.04554595877738, 2.39627597633386, 2.74674301679238, 3.09692650725897,
  -10.2712220944776, -9.92290753816572, -9.57412228338294, -9.22488600047207, 
    -8.87521852517367, -8.5251398520962, -8.1746701280199, -7.82382964504262, 
    -7.4726388335758, -7.12111825519851, -6.76928859537793, 
    -6.41717065606406, -6.06478534816702, -5.71215368392485, 
    -5.35929676917017, -5.00623579550343, -4.65299203238125, 
    -4.29958681912765, -3.94604155687645, -3.59237770045288, 
    -3.23861675020253, -2.88478024377565, -2.5308897478751, 
    -2.17696684997583, -1.82303315002417, -1.4691102521249, 
    -1.11521975622435, -0.761383249797473, -0.407622299547119, 
    -0.0539584431235553, 0.299586819127645, 0.65299203238125, 
    1.00623579550343, 1.35929676917017, 1.71215368392485, 2.06478534816702, 
    2.41717065606406, 2.76928859537793, 3.12111825519851,
  -10.3104526280904, -9.96052962073304, -9.61012812947699, -9.25926813523689, 
    -8.90796978895457, -8.55625340490128, -8.20413945380699, 
    -7.85164855582526, -7.49880147334192, -7.14561910363632, 
    -6.79212247140321, -6.43833272114399, -6.0842711094356, 
    -5.72995899708556, -5.37541784118154, -5.02066918704394, 
    -4.66573466008988, -4.31063595761708, -3.95539484051603, 
    -3.60003312491888, -3.24457267379352, -2.88903538849124, 
    -2.53344320025649, -2.17781806170701, -1.82218193829299, 
    -1.46655679974352, -1.11096461150876, -0.755427326206483, 
    -0.399966875081119, -0.0446051594839685, 0.310635957617082, 
    0.66573466008988, 1.02066918704394, 1.37541784118154, 1.72995899708556, 
    2.0842711094356, 2.43833272114398, 2.79212247140321, 3.14561910363632,
  -10.3501814686258, -9.99863020792764, -9.64659250059007, -9.29408864476818, 
    -8.94113911342926, -8.58776454748223, -8.23398574872706, 
    -7.87982367263292, -7.52529942095383, -7.17043423419068, 
    -6.81524948390831, -6.45976666491649, -6.1040073873235, 
    -5.74799336847125, -5.39174642476052, -5.03528846337529, 
    -4.67864147391481, -4.32182751994225, -3.96486873045871, 
    -3.60778729131134, -3.25060543654442, -2.89334543970212, 
    -2.53602960509168, -2.17868025901598, -1.82131974098402, 
    -1.46397039490832, -1.10665456029789, -0.749394563455581, 
    -0.392212708688666, -0.0351312695412949, 0.321827519942251, 
    0.678641473914813, 1.03528846337529, 1.39174642476052, 1.74799336847125, 
    2.1040073873235, 2.45976666491649, 2.81524948390831, 3.17043423419068,
  -10.3904168913265, -10.0372172628444, -9.683523042678, -9.32935485306493, 
    -8.97473349600169, -8.61967994619524, -8.26421534382698, 
    -7.90836098713838, -7.55213832484746, -7.19556894840521, 
    -6.83867458410108, -6.48147708502679, -6.12399842290749, 
    -5.76626067980946, -5.40828603973349, -5.05009678010311, 
    -4.6917152631568, -4.33316392725328, -3.97446527809912, 
    -3.61564187990769, -3.25671634649874, -2.89771133234766, 
    -2.53864952359353, -2.17955362901525, -1.82044637098475, 
    -1.46135047640647, -1.10228866765234, -0.743283653501258, 
    -0.384358120092313, -0.0255347219008809, 0.333163927253283, 
    0.691715263156799, 1.05009678010311, 1.40828603973349, 1.76626067980946, 
    2.12399842290749, 2.48147708502679, 2.83867458410108, 3.19556894840521,
  -10.431167360405, -10.0762989308818, -9.7209275771652, -9.36507425259594, 
    -9.00876009538868, -8.65200642140011, -8.29483471670181, 
    -7.93726662996736, -7.57932396468325, -7.22102867119308, 
    -6.86240283858456, -6.50346868642891, -6.14424855638207, 
    -5.78476490365741, -5.42504028837928, -5.06509736682705, 
    -4.70495888257916, -4.34464765756663, -3.98418658304563, 
    -3.62359861049857, -3.26290674247337, -2.90213402337018, 
    -2.54130353018542, -2.1804383632223, -1.8195616367777, -1.45869646981458, 
    -1.09786597662982, -0.737093257526632, -0.376401389501426, 
    -0.0158134169543732, 0.344647657566631, 0.704958882579159, 
    1.06509736682705, 1.42504028837928, 1.78476490365741, 2.14424855638207, 
    2.50346868642891, 2.86240283858456, 3.22102867119308,
  -10.4724415343749, -10.1158835449018, -9.75881410592589, -9.40125450909619, 
    -9.04322623622526, -8.68475095186852, -8.32585049570009, 
    -7.96654687469517, -7.60686225512872, -7.24681895440056, 
    -6.88643943269672, -6.52574628449686, -6.16476222993792, 
    -5.80351010604372, -5.44201285783052, -5.08029352929845, 
    -4.71837525431874, -4.35628124742669, -3.99403479453023, 
    -3.63165924354412, -3.2691779949596, -2.90661449235942, 
    -2.54399221288832, -2.18133465768867, -1.81866534231133, 
    -1.45600778711168, -1.09338550764058, -0.730822005040406, 
    -0.368340756455879, -0.00596520546977154, 0.356281247426687, 
    0.718375254318743, 1.08029352929845, 1.44201285783052, 1.80351010604372, 
    2.16476222993792, 2.52574628449685, 2.88643943269671, 3.24681895440056,
  -10.5142482715624, -10.1559796305643, -9.79719081643537, -9.43790346652767, 
    -9.07813941382835, -8.71792067934423, -8.35726946427453, 
    -7.99620814198201, -7.63475924977274, -7.27294548049484, 
    -6.9107896739667, -6.54831480824472, -6.18554399074128, 
    -5.82250044920296, -5.45920752255954, -5.09568865165408, 
    -4.73196736986437, -4.36806729362613, -4.0040121128684, 
    -3.63982558137119, -3.27553150705609, -2.91115374221987, 
    -2.54671617372161, -2.1822427131336, -1.8177572868664, -1.45328382627839, 
    -1.08884625778013, -0.724468492943915, -0.360174418628814, 
    0.00401211286839571, 0.368067293626132, 0.731967369864364, 
    1.09568865165408, 1.45920752255954, 1.82250044920296, 2.18554399074128, 
    2.54831480824472, 2.9107896739667, 3.27294548049484,
  -10.556596635806, -10.1965959118452, -9.83606608709823, -9.47502915221111, 
    -9.11350729912526, -8.75152291326162, -8.38909856548404, 
    -8.02625700385247, -7.66302114517664, -7.29941406638115, 
    -6.9354589956927, -6.57117930366018, -6.2065984940185, -5.84174019440683, 
    -5.47662814695221, -5.11128619872903, -4.74573829210548, 
    -4.38000845498742, -4.01412079097084, -3.64809946941323, 
    -3.28196871543507, -2.91575279986194, -2.54947602911812, 
    -2.1831627350825, -1.8168372649175, -1.45052397088188, -1.08424720013806, 
    -0.718031284564929, -0.351900530586772, 0.0141207909708368, 
    0.380008454987422, 0.745738292105474, 1.11128619872903, 1.47662814695221, 
    1.84174019440683, 2.20659849401849, 2.57117930366018, 2.9354589956927, 
    3.29941406638115,
  -10.5994959023517, -10.2377413167435, -9.87544849276057, -9.5126397821356, 
    -9.1493377437534, -8.78556513562865, -8.42134490665338, 
    -8.05670018812525, -7.69165428506786, -7.32623066735449, 
    -6.96045296064626, -6.59434493715614, -6.22793050625006, 
    -5.86123370489615, -5.49427868797359, -5.12708971845221, 
    -4.75969115745402, -4.392107454208, -4.02436313590938, -3.6564827974946, 
    -3.28849109134319, -2.92041271691788, -2.55227241035414, 
    -2.1840949340103, -1.8159050659897, -1.44772758964587, -1.07958728308212, 
    -0.711508908656812, -0.3435172025054, 0.0243631359093829, 
    0.392107454207996, 0.759691157454015, 1.12708971845221, 1.49427868797359, 
    1.86123370489615, 2.22793050625006, 2.59434493715614, 2.96045296064626, 
    3.32623066735449,
  -10.642955563951, -10.2794249831861, -9.91534681041349, -9.5507437664531, 
    -9.18563878533839, -8.82005500608122, -8.45401576419664, 
    -8.08754458299914, -7.720665164682, -7.35340138119159, -6.9857772649082, 
    -6.61781699914528, -6.24954490847866, -5.88098544891753, 
    -5.51216319792898, -5.14310284432768, -4.77382917804251, 
    -4.40436707977185, -4.03474151053924, -3.66497750116112, 
    -3.2951001416384, -2.92513457048352, -2.55510596399487, 
    -2.18503952549005, -1.81496047450995, -1.44489403600513, 
    -1.07486542951648, -0.704899858361603, -0.335022498838876, 
    0.0347415105392421, 0.404367079771848, 0.773829178042506, 
    1.14310284432768, 1.51216319792898, 1.88098544891753, 2.24954490847866, 
    2.61781699914528, 2.9857772649082, 3.35340138119159,
  -10.6869853371699, -10.3216562651383, -9.95577002509589, -9.58934971516562, 
    -9.22241865295774, -8.85500036711573, -8.48711858861143, 
    -8.11879724180177, -7.75006043525929, -7.38093245238872, 
    -7.01143774184185, -6.64160090774277, -6.27144669973602, 
    -5.90100000286946, -5.53028582732451, -5.15932929800564, 
    -4.78815564400157, -4.41679018793027, -4.04525833518003, 
    -3.67358556305889, -3.30179740986453, -2.92991946388696, 
    -2.55797735235614, -2.18599673034688, -1.81400326965312, 
    -1.44202264764386, -1.07008053611304, -0.698202590135468, 
    -0.32641443694111, 0.0452583351800277, 0.416790187930266, 
    0.78815564400157, 1.15932929800564, 1.5302858273245, 1.90100000286946, 
    2.27144669973602, 2.64160090774277, 3.01143774184185, 3.38093245238872,
  -10.7315951689183, -10.364444738927, -9.99672733600428, -9.62846644401274, 
    -9.25968577279773, -8.89040924950738, -8.52066100965085, 
    -8.15046538790782, -7.77984690870209, -7.40883027655175, 
    -7.03744036620907, -6.66570221260246, -6.29364100059358, 
    -5.92128205456217, -5.54865082783144, -5.17577289194675, 
    -4.80267392582029, -4.42937970475469, -4.05591608935804, 
    -3.68230901436336, -3.30858447736506, -2.93476852748529, 
    -2.56088725398287, -2.18696677481757, -1.81303322518244, 
    -1.43911274601713, -1.06523147251471, -0.691415522634945, 
    -0.317690985636644, 0.0559160893580394, 0.429379704754687, 
    0.802673925820289, 1.17577289194674, 1.54865082783144, 1.92128205456217, 
    2.29364100059358, 2.66570221260246, 3.03744036620907, 3.40883027655175,
  -10.7767952432077, -10.4078002097876, -10.0382281628185, -9.6681029805677, 
    -9.29744877401139, -8.9262898779217, -8.55465084168052, 
    -8.18255641983388, -7.81003156240005, -7.43710140494451, 
    -7.06379125843533, -6.69012659889217, -6.31613305684219, 
    -5.94183640659624, -5.56726255535862, -5.19243753218372, 
    -4.81738747679288, -4.44213862826474, -4.06671731361242, 
    -3.69114993626089, -3.31546296443771, -2.93968291949064, 
    -2.56383636414525, -2.18794989071601, -1.81205010928399, 
    -1.43616363585475, -1.06031708050936, -0.684537035562289, 
    -0.308850063739112, 0.0667173136124194, 0.442138628264735, 
    0.817387476792877, 1.19243753218372, 1.56726255535862, 1.94183640659624, 
    2.31613305684219, 2.69012659889217, 3.06379125843533, 3.43710140494451,
  -10.8225959881466, -10.4517327186416, -10.080282152252, -9.70826857055086, 
    -9.33571649478614, -8.96265067672754, -8.58909608922851, 
    -8.21507791651716, -7.84062154422996, -7.46575254920236, 
    -7.09049668902991, -6.71487989141405, -6.33892824330632, 
    -5.96266797986492, -5.58612547323758, -5.2093272211845, 
    -4.83229983555542, -4.45507003063466, -4.07766461136793, 
    -3.70011046148498, -3.32243453153184, -2.94466382682671, 
    -2.56682539535315, -2.1889463156048, -1.8110536843952, -1.43317460464685, 
    -1.05533617317329, -0.677565468468158, -0.299889538515024, 
    0.0776646113679328, 0.455070030634664, 0.832299835555424, 
    1.2093272211845, 1.58612547323758, 1.96266797986492, 2.33892824330632, 
    2.71487989141405, 3.09049668902991, 3.46575254920236,
  -10.8690080831842, -10.4962525491147, -10.1228991848355, -9.74897268436933, 
    -9.37449798862948, -8.9995002760198, -8.62400495273628, 
    -8.24803764278605, -7.87162417773777, -7.49479058621798, 
    -7.11756308316804, -6.7399680588761, -6.36203206779854, 
    -5.98378181718556, -5.60524415552535, -5.22644606082123, 
    -4.84741462871655, -4.46817706048162, -4.08876065087725, 
    -3.70919277590955, -3.32950088049021, -2.94971246601716, 
    -2.56985507788975, -2.1899562929732, -1.8100437070268, -1.43014492211025, 
    -1.05028753398284, -0.67049911950979, -0.290807224090455, 
    0.0887606508772532, 0.468177060481615, 0.847414628716548, 
    1.22644606082123, 1.60524415552535, 1.98378181718556, 2.36203206779853, 
    2.7399680588761, 3.11756308316804, 3.49479058621798,
  -10.9160424666116, -10.5413702348075, -10.1660893819454, -9.79022502389236, 
    -9.41380253088231, -9.0368475178609, -8.65938583451896, 
    -8.28144355503055, -7.90304696751048, -7.52422256320659, 
    -7.14499702544184, -6.76539721832149, -6.38545017522038, 
    -6.00518308706563, -5.6246232904298, -5.2437982554497, -4.86273557358607, 
    -4.48146294523922, -4.10000816723578, -3.71839912020179, 
    -3.33666375583726, -2.9548300841073, -2.57292616036509, 
    -2.19098007242173, -1.80901992757827, -1.42707383963492, 
    -1.0451699158927, -0.663336244162742, -0.28160087979821, 
    0.100008167235778, 0.48146294523922, 0.862735573586072, 1.2437982554497, 
    1.6246232904298, 2.00518308706563, 2.38545017522038, 2.76539721832149, 
    3.14499702544184, 3.52422256320659,
  -10.9637103433319, -10.5870965668259, -10.2098631130845, -9.83203552947246, 
    -9.4536396254691, -9.07470146275012, -8.69524734494421, 
    -8.31530380708103, -7.93489760474607, -7.55405570295844, 
    -7.17280526478721, -6.79117363972233, -6.40918835181584, 
    -6.02687708760928, -5.64426768386314, -5.26138811510409, 
    -4.87826648100597, -4.4949309936203, -4.11140996447214, 
    -3.72773179153718, -3.34392494611586, -2.9600179596204, 
    -2.57603941029051, -2.19201790985377, -1.80798209014623, 
    -1.42396058970949, -1.0399820403796, -0.656075053884137, 
    -0.272268208462816, 0.111409964472145, 0.494930993620303, 
    0.878266481005972, 1.26138811510409, 1.64426768386314, 2.02687708760928, 
    2.40918835181583, 2.79117363972232, 3.17280526478721, 3.55405570295844,
  -11.0120231929097, -10.6334426015852, -10.2542310034284, -9.87441438722235, 
    -9.49401901189522, -9.11307139633059, -8.73159830883865, 
    -8.34962675630444, -7.96718397302998, -7.58429740928666, 
    -7.20099471959456, -6.81730375074519, -6.43325252958416, 
    -6.04886925057049, -5.66418226312895, -5.27922005881202, 
    -4.89401125828814, -4.50858459817259, -4.12296891771781, 
    -3.7371931453794, -3.35128628527472, -2.96527740355031, 
    -2.57919561467489, -2.19307006767439, -1.80692993232561, 
    -1.42080438532511, -1.03472259644969, -0.648713714725283, 
    -0.262806854620605, 0.122968917717804, 0.508584598172593, 
    0.894011258288135, 1.27922005881202, 1.66418226312895, 2.04886925057049, 
    2.43325252958416, 2.81730375074519, 3.20099471959456, 3.58429740928666,
  -11.0609927779124, -10.6804196688972, -10.2992039416468, -9.91737203655903, 
    -9.53495067250188, -9.15196683634416, -8.76844777213192, 
    -8.38442096992729, -7.99991415432711, -7.6149552726789, 
    -7.22957248301121, -6.84379414169583, -6.45764879085904, 
    -6.07116514555931, -5.68437208074869, -5.29729861803521, 
    -4.9099739122636, -4.52242723793157, -4.13468797545913, 
    -3.74678559732798, -3.35874965410858, -2.97060976039192, 
    -2.58239558064352, -2.19413681499679, -1.80586318500321, 
    -1.41760441935648, -1.02939023960808, -0.64125034589142, 
    -0.25321440267202, 0.134687975459126, 0.522427237931571, 
    0.909973912263596, 1.29729861803521, 1.68437208074869, 2.07116514555931, 
    2.45764879085904, 2.84379414169583, 3.22957248301121, 3.6149552726789,
  -11.1106311525558, -10.7280393803537, -10.3447930880126, -9.96091917802602, 
    -9.57644483998977, -9.19139753984469, -8.80580500874854, 
    -8.41969523159515, -8.03309643519875, -7.64603707616174, 
    -7.25854582844388, -6.87065157065099, -6.48238337306138, 
    -6.09377048440793, -5.70484231843403, -5.31562844024146, 
    -4.92615855244827, -4.53646248117478, -4.14657016187575, 
    -3.7565116250369, -3.36631698175378, -2.97601640921113, 
    -2.58564013608087, -2.19521842785666, -1.80478157214334, 
    -1.41435986391913, -1.02398359078887, -0.633683018246224, 
    -0.243488374963099, 0.146570161875753, 0.536462481174782, 
    0.926158552448273, 1.31562844024146, 1.70484231843403, 2.09377048440793, 
    2.48238337306138, 2.87065157065099, 3.25854582844388, 3.64603707616174,
  -11.1609506716648, -10.7763136380184, -10.3910098828107, -10.0050667814059, 
    -9.61851200522297, -9.23137351068123, -8.8436795277584, 
    -8.45545854817926, -8.06673931325431, -7.67755080138725, 
    -7.28792221527021, -6.8978829687856, -6.50746267363352, 
    -6.11669112570379, -5.72559829121126, -5.33421429261361, 
    -4.94256939433038, -4.55069398828217, -4.15861857926906, 
    -3.76637377020704, -3.37399024724142, -2.98149876475617, 
    -2.58893013029811, -2.1963151894348, -1.8036848105652, -1.41106986970189, 
    -1.01850123524383, -0.626009752758584, -0.233626229792963, 
    0.158618579269058, 0.550693988282166, 0.942569394330378, 
    1.33421429261361, 1.72559829121126, 2.11669112570379, 2.50746267363352, 
    2.8978829687856, 3.28792221527021, 3.67755080138725,
  -11.2119639999661, -10.8252546434401, -10.437866055059, -10.049826094136, 
    -9.6611629253254, -9.27190500726258, -8.88208108079721, 
    -8.49172015684087, -8.1008515038482, -7.70950463495148, -7.3177092947686, 
    -6.92549544590406, -6.53289325516284, -6.13993307949701, 
    -5.74664545170477, -5.35306106590187, -4.959210762785, -4.56512551470718, 
    -4.17083641058478, -3.77637464065605, -3.38177148111097, 
    -2.98705827861213, -2.59226643472661, -2.19742739028842, 
    -1.80257260971158, -1.40773356527339, -1.01294172138787, 
    -0.618228518889035, -0.223625359343951, 0.170836410584777, 
    0.565125514707179, 0.959210762785001, 1.35306106590187, 1.74664545170477, 
    2.13993307949701, 2.53289325516284, 2.92549544590406, 3.3177092947686, 
    3.70950463495147,
  -11.2636841217242, -10.8748749070019, -10.4853736315557, -10.0952086500392, 
    -9.70440863208248, -9.31300255061582, -8.92101966976879, 
    -8.52848953236485, -8.13544194703275, -7.74190697495524, 
    -7.34791491627594, -6.95349629618484, -6.55868185070349, 
    -6.16350251219028, -5.7679893945868, -5.37217377842582, 
    -4.97608709562166, -4.57976091406378, -4.18322692203412, 
    -3.78651691246912, -3.3896627670869, -2.99269644040065, 
    -2.59564994363859, -2.19855532859152, -1.80144467140848, 
    -1.40435005636141, -1.00730355959935, -0.6103372329131, 
    -0.213483087530886, 0.183226922034122, 0.579760914063775, 
    0.976087095621656, 1.37217377842581, 1.7679893945868, 2.16350251219028, 
    2.55868185070349, 2.95349629618484, 3.34791491627594, 3.74190697495524,
  -11.3161243507364, -10.9251872576203, -10.5335449462673, -10.1412262783862, 
    -9.74826044066154, -9.35467693275166, -8.96050555484183, 
    -8.56577639477461, -8.17051981477871, -7.7747664378182, 
    -7.37854713358379, -6.98189300414789, -6.58483536930499, 
    -6.18740575161925, -5.78963586120089, -5.39155758023302, 
    -4.99320294727083, -4.5946041413345, -4.19579346581787, 
    -3.79680333223425, -3.39766624382136, -2.99841477902684, 
    -2.59908157489617, -2.19969931038468, -1.80030068961532, 
    -1.40091842510383, -1.00158522097316, -0.602333756178637, 
    -0.203196667765749, 0.195793465817867, 0.594604141334503, 
    0.993202947270827, 1.39155758023302, 1.78963586120089, 2.18740575161925, 
    2.58483536930499, 2.98189300414789, 3.37854713358379, 3.77476643781819,
  -11.3692983407027, -10.9762048528099, -10.5823926500712, -10.1878911133003, 
    -9.79272995866504, -9.39693922535031, -9.00054926275401, 
    -8.6035907172408, -8.20609451847523, -7.80809186535736, 
    -7.40961421158355, -7.01069325085507, -6.61136090175731, 
    -6.21164929233226, -5.81159074436711, -5.41121775742143, 
    -5.01056299261593, -4.60965925620533, -4.20853948295815, 
    -3.80723671936611, -3.40578410670584, -3.00421486397565, 
    -2.60256227073006, -2.20085964983482, -1.79914035016518, 
    -1.39743772926995, -0.995785136024351, -0.594215893294156, 
    -0.192763280633886, 0.208539482958151, 0.609659256205329, 
    1.01056299261593, 1.41121775742143, 1.81159074436711, 2.21164929233226, 
    2.61136090175731, 3.01069325085507, 3.40961421158355, 3.80809186535736,
  -11.4232200959871, -11.0279411891286, -10.6319297208697, -10.2352156035231, 
    -9.83782909553131, -9.43980078878222, -9.04116159543763, 
    -8.64194273429716, -8.24217571672204, -7.84189233214245, 
    -7.44112463317217, -7.03990492035434, -6.63826572656221, 
    -6.23623980107851, -5.83386009337748, -5.43115973663308, 
    -5.02817203097741, -4.62493042653305, -4.22146850624302, 
    -3.8178199685224, -3.41401860975512, -3.01009830665997, 
    -2.60609299854944, -2.2020366695053, -1.7979633304947, -1.39390700145056, 
    -0.989901693340028, -0.585981390244877, -0.182180031477602, 
    0.22146850624302, 0.624930426533046, 1.02817203097741, 1.43115973663308, 
    1.83386009337748, 2.23623980107851, 2.63826572656221, 3.03990492035434, 
    3.44112463317217, 3.84189233214245,
  -11.4779039827867, -11.0804101130221, -10.6821694740909, -10.2832125225558, 
    -9.88357007229861, -9.48327328147863, -9.08235363898089, 
    -8.68084295037736, -8.27877332342718, -7.87617715314035, 
    -7.47308710643013, -7.06953610637869, -6.66555731614141, 
    -6.26118412251436, -5.85645011919016, -5.45138908972704, 
    -5.04603499025606, -4.64042193195145, -4.23458416328895, 
    -3.82855605211717, -3.42237206756684, -3.01606676182288, 
    -2.60967475178431, -2.20323070063685, -1.79676929936315, 
    -1.39032524821569, -0.983933238177125, -0.577627932433165, 
    -0.171443947882831, 0.234584163288947, 0.640421931951449, 
    1.04603499025606, 1.45138908972704, 1.85645011919016, 2.26118412251436, 
    2.66555731614141, 3.06953610637869, 3.47308710643012, 3.87617715314035,
  -11.5333647407262, -11.1336258320837, -10.7331255735949, -10.3318949791922, 
    -9.92996543174863, -9.527368669668, -9.12413677294049, -8.72030214868767, 
    -8.31589751622423, -7.91095589166232, -7.50551057208454, 
    -7.09959511931187, -6.69324334329251, -6.28648928513789, 
    -5.87936719983203, -5.47191153864015, -5.06415693124302, 
    -4.6561381676228, -4.24789017972691, -3.83944802293568, 
    -3.43084685736024, -3.02212192899656, -2.61330855076194, 
    -2.20444208343995, -1.79555791656005, -1.38669144923806, 
    -0.977878071003439, -0.569153142639765, -0.160551977064324, 
    0.247890179726906, 0.6561381676228, 1.06415693124302, 1.47191153864015, 
    1.87936719983203, 2.28648928513789, 2.6932433432925, 3.09959511931187, 
    3.50551057208454, 3.91095589166232,
  -11.589617494899, -11.1876029267477, -10.7848120430015, -10.3812764284626, 
    -9.9770280489468, -9.57209923749472, -9.16652268002128, 
    -8.76033140043058, -8.35355874522382, -7.94623836762767, 
    -7.5384042112704, -7.13009049343321, -6.72133168790423, 
    -6.31216250746245, -5.90261788601917, -5.49273296044418, 
    -5.08254305210431, -4.67208364814145, -4.26139038251782, 
    -3.85049901685548, -3.43944542109792, -3.02826555402072, 
    -2.61699544361902, -2.20567116739903, -1.79432883260097, 
    -1.38300455638098, -0.971734445979285, -0.560554578902085, 
    -0.149500983144521, 0.261390382517814, 0.672083648141453, 
    1.08254305210431, 1.49273296044418, 1.90261788601916, 2.31216250746245, 
    2.72133168790423, 3.13009049343321, 3.5384042112704, 3.94623836762767,
  -11.6466777683717, -11.2423563624383, -10.8372432774614, -10.4313706830064, 
    -10.0247711421974, -9.61747759753784, -9.20952335614008, 
    -8.80094207439598, -8.39176774211491, -7.98203466615899, 
    -7.57177745360397, -7.16103099445463, -6.7498304439433, 
    -6.33821120444043, -5.92620890700573, -5.51385939260887, 
    -5.10119869304827, -4.68826301159688, -4.27508870340356, 
    -3.86171225567894, -3.44817026769444, -3.0344994306231, 
    -2.62073650725122, -2.20691831158922, -1.79308168841078, 
    -1.37926349274878, -0.965500569376899, -0.551829732305564, 
    -0.138287744321057, 0.275088703403558, 0.68826301159688, 
    1.10119869304827, 1.51385939260887, 1.92620890700573, 2.33821120444043, 
    2.7498304439433, 3.16103099445463, 3.57177745360397, 3.98203466615899,
  -11.704561495175, -11.2979015021913, -10.8904340558877, -10.4821919248927, 
    -10.0732082844328, -9.66351670174817, -9.25315112089137, 
    -8.84214584693667, -8.43053552963219, -8.01835514652411, 
    -7.60563998558315, -7.19242562736373, -6.77874792672573, 
    -6.3646429941492, -5.95014717667198, -5.53529703848063, 
    -5.12012934118455, -4.70468102380373, -4.28898918250006, 
    -3.87309105008246, -3.45702397531606, -3.04082540206539, 
    -2.62453284830193, -2.20818388500611, -1.79181611499389, 
    -1.37546715169807, -0.959174597934615, -0.542976024683939, 
    -0.126908949917538, 0.288989182500055, 0.704681023803729, 
    1.12012934118455, 1.53529703848062, 1.95014717667198, 2.3646429941492, 
    2.77874792672573, 3.19242562736373, 3.60563998558315, 4.01835514652411,
  -11.7632850338022, -11.3542541197723, -10.9443995536712, -10.533754717911, 
    -10.1223534150559, -9.71022985282315, -9.29741862843367, 
    -8.88395471234645, -8.46987343140692, -8.05521045144154, 
    -7.64000175933011, -7.22428364458744, -6.80809268048607, 
    -6.39146570475173, -5.97443979986303, -5.55705227298728, 
    -5.13934063558387, -4.72134258270699, -4.30309597203926, 
    -3.88463880268806, -3.46600919377599, -3.04724536285737, 
    -2.62838560419217, -2.20946826690931, -1.79053173309069, 
    -1.37161439580783, -0.952754637142635, -0.533990806224006, 
    -0.11536119731194, 0.303095972039261, 0.721342582706984, 
    1.13934063558387, 1.55705227298728, 1.97443979986303, 2.39146570475173, 
    2.80809268048607, 3.22428364458744, 3.64000175933011, 4.05521045144154,
  -11.8228651812381, -11.4114304133135, -10.9991553559011, -10.5860740203507, 
    -10.1722208522589, -9.75763071604006, -9.3423388788163, 
    -8.92638099365967, -8.50979308221917, -8.09261151676635, 
    -7.67487300169265, -7.25661455449158, -6.83787348625905, 
    -6.41868738174513, -5.99909407899034, -5.5791316485798, 
    -5.15883837254848, -4.73825272297074, -4.31741334026735, 
    -3.89635901126333, -3.47512864702979, -3.05376126054293, 
    -2.63229594419356, -2.2107718471803, -1.7892281528197, -1.36770405580644, 
    -0.946238739457075, -0.52487135297021, -0.103640988736668, 
    0.317413340267346, 0.738252722970738, 1.15883837254848, 1.57913164857979, 
    1.99909407899034, 2.41868738174513, 2.83787348625905, 3.25661455449158, 
    3.67487300169265, 4.09261151676635,
  -11.8833191875431, -11.4694470194926, -11.0547174711133, -10.6391651982963, 
    -10.222825305838, -9.80573333156889, -9.38792522976725, 
    -8.96943735389218, -8.55030643867084, -8.13056958157496, 
    -7.71026422372155, -7.28942813023258, -6.86809937008857, 
    -6.44631629551106, -6.02411752090878, -5.60154190142249, 
    -5.17862851110332, -4.75541662075953, -4.3319456755067, 
    -3.90825527205601, -3.48438513577584, -3.06037509756126, 
    -2.63626507054653, -2.21209502669548, -1.78790497330452, 
    -1.36373492945347, -0.939624902438742, -0.51561486422416, 
    -0.0917447279439912, 0.331945675506695, 0.755416620759534, 
    1.17862851110332, 1.60154190142249, 2.02411752090878, 2.44631629551105, 
    2.86809937008857, 3.28942813023258, 3.71026422372155, 4.13056958157496,
  -11.9446647710174, -11.5283210282795, -11.1111023455931, -10.6930440394583, 
    -10.2741818905294, -9.85455212728789, -9.43419140896436, 
    -9.01313680774492, -8.59142579029939, -8.16909619866781, 
    -7.74618623054194, -7.3227344189784, -6.89877961158009, -6.4743609491827, 
    -6.04951784408274, -5.62428995784402, -5.19871717871897, 
    -4.7728395987218, -4.34669749038982, -3.92033128326982, 
    -3.49378154016616, -3.06708893318707, -2.64029421962607, 
    -2.21343821771492, -1.78656178228508, -1.35970578037393, 
    -0.932911066812927, -0.506218459833841, -0.0796687167301795, 
    0.346697490389816, 0.772839598721802, 1.19871717871897, 1.62428995784402, 
    2.04951784408274, 2.4743609491827, 2.89877961158009, 3.3227344189784, 
    3.74618623054194, 4.16909619866781,
  -12.0069201339725, -11.5880699982758, -11.1683268782555, -10.7477267675679, 
    -10.3263061398906, -9.90410193212539, -9.48115152681256, 
    -9.05749273379225, -8.63316377115382, -8.20820324551046, 
    -7.78265013163804, -7.35654375151665, -6.92992375281321, 
    -6.50283008684404, -6.07530298605556, -5.64738294106189, 
    -5.21911067727776, -4.79052713118539, -4.36167342627371, 
    -3.93259084868867, -3.50332082263294, -3.07390488555373, 
    -2.6443846631572, -2.21480184428792, -1.78519815571208, -1.3556153368428, 
    -0.92609511444627, -0.496679177367065, -0.0674091513113325, 
    0.36167342627371, 0.790527131185385, 1.21911067727776, 1.64738294106189, 
    2.07530298605556, 2.50283008684404, 2.92992375281321, 3.35654375151664, 
    3.78265013163804, 4.20820324551045,
  -12.070103979138, -11.6487119726777, -11.2264084361333, -10.8032300573612, 
    -10.3792140207527, -9.95439798995343, -9.5288200897519, 
    -9.10251888717863, -8.67553337185514, -8.24790293563419, 
    -7.81966735157143, -7.39086675226909, -6.96154160763217, 
    -6.53173270207764, -6.10148111123723, -5.67082817819428, 
    -5.23981548929516, -4.80848484957577, -4.37687825784371, 
    -3.94503788145654, -3.51300603083667, -3.08082513376345, 
    -2.64853770948295, -2.21618634267585, -1.78381365732415, 
    -1.35146229051705, -0.919174866236546, -0.48699396916333, 
    -0.0549621185434572, 0.376878257843714, 0.808484849575768, 
    1.23981548929515, 1.67082817819428, 2.10148111123723, 2.53173270207764, 
    2.96154160763217, 3.39086675226909, 3.81966735157143, 4.24790293563418,
  -12.1342355267336, -11.7102654958874, -11.2853648704987, -10.8595710501805, 
    -10.4329219482722, -10.0054559740595, -9.57721201412183, 
    -9.14822941284821, -8.71854795216523, -8.28820783051903, 
    -7.85724964115423, -7.42571434973251, -6.99364327133317, 
    -6.56107804687848, -6.12806061902643, -5.69463320757339, 
    -5.26083828440931, -4.8267185480682, -4.39231689791638, 
    -3.95767640802106, -3.52284030074205, -3.08785192008905, 
    -2.65275470488719, -2.21759216179346, -1.78240783820654, 
    -1.34724529511281, -0.912148079910951, -0.477159699257949, 
    -0.0423235919789379, 0.392316897916384, 0.826718548068204, 
    1.2608382844093, 1.69463320757339, 2.12806061902643, 2.56107804687848, 
    2.99364327133316, 3.42571434973251, 3.85724964115423, 4.28820783051902,
  -12.1993345322379, -11.7727496308086, -11.3452145336514, -10.9167673702236, 
    -10.487446801609, -10.0572920022249, -9.62634264060909, 
    -9.19463885933374, -8.76222125408908, -8.32913085198284, 
    -7.89540908909996, -7.46109778736727, -7.02623913076819, 
    -6.59087564095217, -6.15505015228367, -5.71880578637566, 
    -5.28218592615226, -4.84523418948561, -4.40799440245151, 
    -3.97051057224892, -3.53282685982804, -3.09498755227176, 
    -2.65703703497538, -2.21901976366946, -1.78098023633054, 
    -1.34296296502462, -0.905012447728242, -0.467173140171956, 
    -0.0294894277510777, 0.407994402451507, 0.845234189485611, 
    1.28218592615226, 1.71880578637565, 2.15505015228367, 2.59087564095217, 
    3.02623913076819, 3.46109778736727, 3.89540908909996, 4.32913085198284,
  -12.2654213048853, -11.8361839768544, -11.4059762964037, -10.9748371414709, 
    -10.542805940264, -10.1099226524386, -9.67622774930778, 
    -9.24176219313222, -8.80656741553677, -8.37068529510182, 
    -7.93415813417573, -7.49702863495608, -7.05933987488657, 
    -6.62113528141696, -6.18245860617323, -5.74335389858492, 
    -5.30386547901725, -4.86403791145476, -4.42391597578396, 
    -3.98354463972209, -3.54296903043911, -3.10223440592021, 
    -2.66138612611596, -2.22046962392733, -1.77953037607267, 
    -1.33861387388404, -0.897765594079794, -0.457030969560894, 
    -0.0164553602779117, 0.423915975783961, 0.86403791145476, 
    1.30386547901725, 1.74335389858492, 2.18245860617322, 2.62113528141696, 
    3.05933987488657, 3.49702863495608, 3.93415813417573, 4.37068529510182,
  -12.3325167269287, -11.9005886887045, -11.4676695662959, -11.0337990053248, 
    -10.599017221106, -10.163364979279, -9.72688357542193, -9.28961481369649, 
    -8.85160098457344, -8.41288484168897, -7.97350957788124, 
    -7.53351880045672, -7.09295650573622, -6.65186705293018, 
    -6.21029513739293, -5.76828576330557, -5.32588421583718, 
    -4.88313603283407, -4.44008697608672, -3.99678300222404, 
    -3.5532702332848, -3.10959492701567, -2.66580344694581, 
    -2.22194223228748, -1.77805776771252, -1.33419655305419, 
    -0.890405072984334, -0.446729766715203, -0.00321699777595758, 
    0.440086976086718, 0.883136032834071, 1.32588421583718, 1.76828576330557, 
    2.21029513739293, 2.65186705293018, 3.09295650573622, 3.53351880045672, 
    3.97350957788124, 4.41288484168897,
  -12.4006422737013, -11.9659844958466, -11.5303143065788, -11.0936721389949, 
    -10.6560990161236, -10.2176365309956, -9.77832682564251, 
    -9.33821256907373, -8.89733693428639, -8.45574357435891, 
    -8.01347659768122, -7.57058054237387, -7.12710034994831, 
    -6.68308133826069, -6.23856917381156, -5.79360984344368, 
    -5.34824962549043, -4.90253506042705, -4.456512921077, -4.01023018242595, 
    -3.5637339910955, -3.11707163452915, -2.67029050994277, 
    -2.22343809309188, -1.77656190690812, -1.32970949005723, 
    -0.882928365470851, -0.436266008904503, 0.0102301824259485, 
    0.456512921077001, 0.902535060427047, 1.34824962549043, 1.79360984344368, 
    2.23856917381156, 2.68308133826069, 3.12710034994831, 3.57058054237387, 
    4.01347659768122, 4.45574357435891,
  -12.4698200345189, -12.032392722941, -11.5939310560001, -11.1544762746665, 
    -10.7140702309367, -10.2727553673263, -9.83057469523287, 
    -9.38757177222333, -8.94379067830114, -8.49927599120867, 
    -8.05407276081961, -7.60822648267676, -7.16178307073012, 
    -6.71478882933073, -6.26729042453506, -5.81933485477538, 
    -5.37096942095112, -4.92224169599629, -4.47319949397832, 
    -4.02389083878324, -3.57436393244245, -3.12466712315623, 
    -2.67484887306912, -2.22495772585223, -1.77504227414778, 
    -1.32515112693088, -0.875332876843769, -0.425636067557554, 
    0.0238908387832375, 0.473199493978319, 0.922241695996286, 
    1.37096942095111, 1.81933485477538, 2.26729042453506, 2.71478882933073, 
    3.16178307073012, 3.60822648267676, 4.05407276081961, 4.49927599120867,
  -12.5400727344615, -12.0998353110477, -11.6585409494342, -11.216231719491, 
    -10.7729503241066, -10.328740078086, -9.88364488585808, 
    -9.43770921804868, -8.99097808697895, -8.54349702114615, 
    -8.09531203874544, -7.64646962029068, -7.19701668039243, 
    -6.74700053875116, -6.29646889042395, -5.84546977542262, 
    -5.39405154770167, -4.94226284359386, -4.49015254975182, 
    -4.03776977065366, -3.58516379573075, -3.1323840661758, 
    -2.67948014148939, -2.22650166582304, -1.77349833417696, 
    -1.32051985851061, -0.867615933824202, -0.414836204269249, 
    0.0377697706536641, 0.490152549751822, 0.942262843593857, 
    1.39405154770167, 1.84546977542262, 2.29646889042394, 2.74700053875116, 
    3.19701668039243, 3.64646962029068, 4.09531203874543, 4.54349702114615,
  -12.6114237570777, -12.1683348397586, -11.724165739397, -11.2789593764394, 
    -10.8327593272841, -10.3856098025678, -9.93755562419635, 
    -9.48864220117936, -9.0389155043313, -8.58842203989972, 
    -8.13720882218208, -7.68532334519246, -7.23281355343942, 
    -6.77972781187636, -6.32611487508564, -5.8720238557578, -5.4175041925271, 
    -4.9626056172248, -4.5073781216113, -4.05187192364866, -3.59613743337458, 
    -3.14022521843934, -2.6841859693668, -2.22807046460093, 
    -1.77192953539907, -1.3158140306332, -0.859774781560662, 
    -0.40386256662542, 0.0518719236486579, 0.507378121611304, 
    0.962605617224802, 1.4175041925271, 1.8720238557578, 2.32611487508564, 
    2.77972781187636, 3.23281355343942, 3.68532334519246, 4.13720882218208, 
    4.58842203989972 ;

 projection_x_coordinate = -187500, -162500, -137500, -112500, -87500, 
    -62500, -37500, -12500, 12500, 37500, 62500, 87500, 112500, 137500, 
    162500, 187500, 212500, 237500, 262500, 287500, 312500, 337500, 362500, 
    387500, 412500, 437500, 462500, 487500, 512500, 537500, 562500, 587500, 
    612500, 637500, 662500, 687500, 712500, 737500, 762500 ;

 projection_x_coordinate_bnds =
  -200000, -175000,
  -175000, -150000,
  -150000, -125000,
  -125000, -100000,
  -100000, -75000,
  -75000, -50000,
  -50000, -25000,
  -25000, 0,
  0, 25000,
  25000, 50000,
  50000, 75000,
  75000, 100000,
  100000, 125000,
  125000, 150000,
  150000, 175000,
  175000, 200000,
  200000, 225000,
  225000, 250000,
  250000, 275000,
  275000, 300000,
  300000, 325000,
  325000, 350000,
  350000, 375000,
  375000, 400000,
  400000, 425000,
  425000, 450000,
  450000, 475000,
  475000, 500000,
  500000, 525000,
  525000, 550000,
  550000, 575000,
  575000, 600000,
  600000, 625000,
  625000, 650000,
  650000, 675000,
  675000, 700000,
  700000, 725000,
  725000, 750000,
  750000, 775000 ;

 projection_y_coordinate = -87500, -62500, -37500, -12500, 12500, 37500, 
    62500, 87500, 112500, 137500, 162500, 187500, 212500, 237500, 262500, 
    287500, 312500, 337500, 362500, 387500, 412500, 437500, 462500, 487500, 
    512500, 537500, 562500, 587500, 612500, 637500, 662500, 687500, 712500, 
    737500, 762500, 787500, 812500, 837500, 862500, 887500, 912500, 937500, 
    962500, 987500, 1012500, 1037500, 1062500, 1087500, 1112500, 1137500, 
    1162500, 1187500 ;

 projection_y_coordinate_bnds =
  -100000, -75000,
  -75000, -50000,
  -50000, -25000,
  -25000, 0,
  0, 25000,
  25000, 50000,
  50000, 75000,
  75000, 100000,
  100000, 125000,
  125000, 150000,
  150000, 175000,
  175000, 200000,
  200000, 225000,
  225000, 250000,
  250000, 275000,
  275000, 300000,
  300000, 325000,
  325000, 350000,
  350000, 375000,
  375000, 400000,
  400000, 425000,
  425000, 450000,
  450000, 475000,
  475000, 500000,
  500000, 525000,
  525000, 550000,
  550000, 575000,
  575000, 600000,
  600000, 625000,
  625000, 650000,
  650000, 675000,
  675000, 700000,
  700000, 725000,
  725000, 750000,
  750000, 775000,
  775000, 800000,
  800000, 825000,
  825000, 850000,
  850000, 875000,
  875000, 900000,
  900000, 925000,
  925000, 950000,
  950000, 975000,
  975000, 1000000,
  1000000, 1025000,
  1025000, 1050000,
  1050000, 1075000,
  1075000, 1100000,
  1100000, 1125000,
  1125000, 1150000,
  1150000, 1175000,
  1175000, 1200000 ;

 time = 1586976, 1587720, 1588392, 1589136, 1589856, 1590600, 1591320, 
    1592064, 1592808, 1593528, 1594272, 1594992 ;

 season_year = 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;
}
