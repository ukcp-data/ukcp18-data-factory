netcdf ukcp18-land-gcm-uk-river-mon {
dimensions:
	ensemble_member = 1 ;
	region = 26 ;
	strlen = 21 ;
	time = 12 ;
	bnds = 2 ;
variables:
	float ensemble_member(ensemble_member) ;
		ensemble_member:units = "" ;
		ensemble_member:long_name = "Ensemble member" ;
	float example_var(ensemble_member, time, region) ;
		example_var:_FillValue = 1.e+20f ;
		example_var:standard_name = "air_temperature" ;
		example_var:long_name = "Monthly mean air temperature" ;
		example_var:units = "degC" ;
		example_var:cell_methods = "time: mid_range within days time: mean over days" ;
		example_var:coordinates = "geo_region" ;
	char geo_region(region, strlen) ;
		geo_region:standard_name = "region" ;
		geo_region:long_name = "River basin" ;
	double time(time) ;
		time:axis = "T" ;
		time:units = "hours since 1851-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "standard" ;

// global attributes:
		:comment = "These data are part of the test suite for the data-factory." ;
		:references = "" ;
		:short_name = "temp data" ;
		:source = "a project" ;
		:title = "Great data at your service" ;
		:Conventions = "CF-1.5" ;
data:

 ensemble_member = 1 ;

 example_var =
  7.03, 6.89, 6.17, 5.3, 4.54, 4.92, 5.84, 5.18, 4.15, 4.32, 5.04, 4.7, 4.68, 
    1.42, 3.72, 3.69, 4.14, 4.19, 4.44, 2.85, 3.88, 4.15, 3.74, 4.37, 3.91, 
    3.87,
  2.95, 4.62, 3.22, 4.45, 3.99, 4.3, 4.56, 2.43, 4.29, 3.88, 4.76, 3.25, 
    3.91, 4.22, 4.6, 5.17, 2.7, 2.37, 4.73, 4.35, 3.73, 2.81, 3.49, 1.85, 
    7.94, 8.04,
  7.53, 7.16, 6.23, 7.01, 6.51, 6.44, 6.6, 4.08, 6.64, 6.32, 6.52, 5.27, 
    6.22, 5.97, 6.51, 6.75, 4.59, 4.17, 6.58, 6.19, 5.49, 4.39, 4.44, 4.93, 
    6.4, 4.68,
  2.98, 5.71, 3.83, 3.91, 5.97, 4.21, 2.1, 3.47, 3.48, 6.07, 2.78, 2.15, 1.7, 
    1.87, 5.48, 4.5, 3.31, 9.07, 9.4, 8.88, 8.86, 8.04, 8.93, 9.72, 9.27, 8.26,
  8.56, 9.38, 8.85, 8.16, 4.47, 7.59, 7.77, 8.44, 8.61, 9.02, 6.33, 8.06, 
    8.38, 8.19, 8.95, 8.36, 8.5, 5.98, 8.72, 7.41, 8.89, 8.51, 8.45, 8.68, 
    6.25, 8.69,
  8.23, 8.71, 7.38, 8.23, 7.77, 8.24, 8.42, 6.58, 6.16, 8.23, 7.92, 7.47, 
    6.42, 6.65, 6.77, 8.24, 6.82, 5.03, 7.49, 5.98, 6.21, 7.84, 6.13, 4.42, 
    5.71, 5.73,
  7.86, 4.93, 4.24, 3.79, 4.02, 7.36, 6.39, 5.36, 11.61, 12.26, 11.71, 11.88, 
    11.25, 12.2, 13.07, 12.5, 11.45, 11.76, 12.71, 12.13, 11.12, 7.62, 10.36, 
    11.08, 11.61, 11.82,
  12.24, 9.33, 11.14, 11.62, 11.31, 12.1, 11.59, 11.67, 8.91, 11.79, 10.57, 
    12.02, 11.62, 11.51, 11.85, 9.66, 11.73, 11.21, 12, 10.52, 11.27, 10.46, 
    10.89, 11, 9.53, 9.05,
  10.93, 10.43, 10.32, 9.25, 9.56, 9.45, 11.02, 9.7, 7.83, 9.97, 8.95, 9.23, 
    10.43, 8.86, 7.42, 8.62, 8.43, 10.45, 7.79, 6.97, 6.48, 6.88, 9.81, 9.07, 
    7.94, 13.98,
  14.83, 14.21, 14.65, 13.97, 15, 15.93, 15.4, 14.34, 14.68, 15.68, 15.1, 
    13.64, 10.02, 13.26, 14.01, 14.58, 14.81, 15.23, 11.88, 13.96, 14.45, 
    14.26, 15.05, 14.5, 14.63, 11.41,
  14.49, 13.29, 14.95, 14.53, 14.34, 14.41, 12.19, 14.7, 14.2, 14.5, 13.23, 
    14.14, 13, 13.57, 13.58, 12.15, 11.89, 13.68, 13.01, 12.85, 11.87, 12.14, 
    12.2, 13.38, 12.23, 10.52,
  12.64, 11.35, 11.67, 13.08, 10.91, 9.68, 11.29, 11.1, 12.53, 10.26, 9.7, 
    9.15, 9.17, 12.48, 11.18, 10.36, 15.97, 16.87, 16.22, 16.66, 16.05, 
    17.13, 18.15, 17.36, 16.52, 16.98 ;

 geo_region =
  "argyll",
  "tay",
  "orkney_and_shetlands",
  "north_east_scotland",
  "anglian",
  "channel_islands",
  "isle_of_man",
  "clyde",
  "north_western_ireland",
  "south_east_england",
  "west_highland",
  "tweed",
  "forth",
  "north_eastern_ireland",
  "northumbria",
  "humber",
  "north_highland",
  "south_west_england",
  "north_west_england",
  "solway",
  "west_wales",
  "republic_of_ireland",
  "neagh_bann",
  "thames",
  "severn",
  "dee" ;

 time = 1586976, 1587720, 1588392, 1589136, 1589856, 1590600, 1591320, 
    1592064, 1592808, 1593528, 1594272, 1594992 ;
}
