netcdf ukcp18-land-gcm-uk-60km-mon {
dimensions:
	ensemble_member = 1 ;
	time = 12 ;
	bnds = 2 ;
	projection_y_coordinate = 25 ;
	projection_x_coordinate = 15 ;
variables:
	float ensemble_member(ensemble_member) ;
		ensemble_member:units = "" ;
		ensemble_member:long_name = "Ensemble member" ;
	float example_var(ensemble_member, time, projection_y_coordinate, projection_x_coordinate) ;
		example_var:_FillValue = 1.e+20f ;
		example_var:standard_name = "air_temperature" ;
		example_var:long_name = "Monthly mean air temperature" ;
		example_var:units = "degC" ;
		example_var:cell_methods = "time: mid_range within days time: mean over days" ;
		example_var:coordinates = "latitude longitude" ;
		example_var:grid_mapping = "transverse_mercator" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	double latitude(projection_y_coordinate, projection_x_coordinate) ;
		latitude:units = "degree_north" ;
		latitude:standard_name = "latitude" ;
	double longitude(projection_y_coordinate, projection_x_coordinate) ;
		longitude:units = "degree_east" ;
		longitude:standard_name = "longitude" ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	double time(time) ;
		time:axis = "T" ;
		time:units = "hours since 1851-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "standard" ;
	int season_year(time) ;
		season_year:units = "1" ;
		season_year:long_name = "season_year" ;

// global attributes:
		:comment = "These data are part of the test suite for the data-factory." ;
		:references = "" ;
		:short_name = "temp data" ;
		:source = "a project" ;
		:title = "Great data at your service" ;
		:Conventions = "CF-1.5" ;
		:history = "Fri Oct 13 05:39:26 2017: ncks -d projection_x_coordinate,,,12 -d projection_y_coordinate,,,12 -v example_var osgb_5km.nc osgb_60km.nc" ;
		:NCO = "\"4.5.5\"" ;
data:

 ensemble_member = 1 ;

 example_var =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 7.03, _, 6.89, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 6.17, 5.3, 4.54, 4.92, 5.84, _, _, _,
  _, _, _, _, _, _, _, _, _, 5.18, 4.15, 4.32, 5.04, 4.7, _,
  _, _, _, _, _, _, _, 4.68, 1.42, 3.72, 3.69, 4.14, 4.19, 4.44, _,
  _, _, _, _, _, _, _, _, 2.85, 3.88, 4.15, 3.74, 4.37, 3.91, 3.87,
  _, _, _, _, _, _, _, _, 2.95, 4.62, 3.22, 4.45, 3.99, 4.3, _,
  _, _, _, _, _, _, _, _, _, 4.56, 2.43, 4.29, 3.88, _, _,
  _, _, _, _, _, _, _, _, _, 4.76, 3.25, 3.91, _, _, _,
  _, _, _, _, 4.22, 4.6, 5.17, _, _, 2.7, 2.37, 4.73, _, _, _,
  _, _, _, _, _, 4.35, _, 3.73, 2.81, 2.58, 3.02, _, _, _, _,
  _, _, _, _, _, _, _, 5.31, 2.75, 1.37, 3.72, _, _, _, _,
  _, _, _, _, _, _, _, 2.68, 2.27, 4.14, _, _, _, _, _,
  _, _, _, _, _, _, 3.24, 1.19, 1.55, 1.66, _, _, _, _, _,
  _, _, _, _, _, _, 4.71, 1.27, 0.53, 0.32, _, _, _, _, _,
  _, _, _, _, _, _, _, 0.8, 3.51, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 3.37, 1.85, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 6.76, _, 6.61, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 5.94, 5.23, 4.32, 4.93, 5.68, _, _, _,
  _, _, _, _, _, _, _, _, _, 5.27, 4.13, 4.35, 5.04, 4.57, _,
  _, _, _, _, _, _, _, 4.68, 0.96, 3.61, 3.57, 4.22, 4.17, 4.49, _,
  _, _, _, _, _, _, _, _, 2.62, 3.89, 4.13, 3.79, 4.47, 3.97, 3.96,
  _, _, _, _, _, _, _, _, 2.64, 4.7, 3.27, 4.58, 4.22, 4.36, _,
  _, _, _, _, _, _, _, _, _, 4.64, 2.31, 4.44, 4.17, _, _,
  _, _, _, _, _, _, _, _, _, 4.8, 3.32, 4.16, _, _, _,
  _, _, _, _, 4.33, 4.8, 5.27, _, _, 2.8, 2.38, 4.98, _, _, _,
  _, _, _, _, _, 4.54, _, 3.85, 2.88, 2.79, 3.25, _, _, _, _,
  _, _, _, _, _, _, _, 5.23, 2.98, 1.37, 4.09, _, _, _, _,
  _, _, _, _, _, _, _, 2.73, 2.44, 4.44, _, _, _, _, _,
  _, _, _, _, _, _, 3.11, 1.05, 1.76, 1.94, _, _, _, _, _,
  _, _, _, _, _, _, 4.8, 1.31, 0.6, 0.26, _, _, _, _, _,
  _, _, _, _, _, _, _, 0.68, 3.71, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 3.49, 1.85, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 7.94, _, 8.04, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 7.53, 7.16, 6.23, 7.01, 7.66, _, _, _,
  _, _, _, _, _, _, _, _, _, 7.4, 6.29, 6.62, 7.31, 6.88, _,
  _, _, _, _, _, _, _, 6.42, 2.48, 5.5, 5.72, 6.47, 6.56, 6.88, _,
  _, _, _, _, _, _, _, _, 4.54, 6.09, 6.32, 6.15, 6.92, 6.26, 6.32,
  _, _, _, _, _, _, _, _, 4.22, 6.86, 5.4, 6.85, 6.51, 6.44, _,
  _, _, _, _, _, _, _, _, _, 6.6, 4.08, 6.64, 6.32, _, _,
  _, _, _, _, _, _, _, _, _, 6.52, 5.27, 6.22, _, _, _,
  _, _, _, _, 5.97, 6.51, 6.75, _, _, 4.59, 4.17, 6.58, _, _, _,
  _, _, _, _, _, 6.19, _, 5.49, 4.39, 4.44, 4.93, _, _, _, _,
  _, _, _, _, _, _, _, 6.4, 4.68, 2.98, 5.71, _, _, _, _,
  _, _, _, _, _, _, _, 3.83, 3.91, 5.97, _, _, _, _, _,
  _, _, _, _, _, _, 4.21, 2.1, 3.47, 3.48, _, _, _, _, _,
  _, _, _, _, _, _, 6.07, 2.78, 2.15, 1.7, _, _, _, _, _,
  _, _, _, _, _, _, _, 1.87, 5.48, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 4.5, 3.31, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 9.07, _, 9.4, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 8.88, 8.86, 8.04, 8.93, 9.72, _, _, _,
  _, _, _, _, _, _, _, _, _, 9.27, 8.26, 8.56, 9.38, 8.85, _,
  _, _, _, _, _, _, _, 8.16, 4.47, 7.59, 7.77, 8.44, 8.61, 9.02, _,
  _, _, _, _, _, _, _, _, 6.33, 8.06, 8.38, 8.19, 8.95, 8.36, 8.5,
  _, _, _, _, _, _, _, _, 5.98, 8.72, 7.41, 8.89, 8.51, 8.45, _,
  _, _, _, _, _, _, _, _, _, 8.68, 6.25, 8.69, 8.23, _, _,
  _, _, _, _, _, _, _, _, _, 8.71, 7.38, 8.23, _, _, _,
  _, _, _, _, 7.77, 8.24, 8.42, _, _, 6.58, 6.16, 8.23, _, _, _,
  _, _, _, _, _, 7.92, _, 7.47, 6.42, 6.65, 6.77, _, _, _, _,
  _, _, _, _, _, _, _, 8.24, 6.82, 5.03, 7.49, _, _, _, _,
  _, _, _, _, _, _, _, 5.98, 6.21, 7.84, _, _, _, _, _,
  _, _, _, _, _, _, 6.13, 4.42, 5.71, 5.73, _, _, _, _, _,
  _, _, _, _, _, _, 7.86, 4.93, 4.24, 3.79, _, _, _, _, _,
  _, _, _, _, _, _, _, 4.02, 7.36, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 6.39, 5.36, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 11.61, _, 12.26, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 11.71, 11.88, 11.25, 12.2, 13.07, _, _, _,
  _, _, _, _, _, _, _, _, _, 12.5, 11.45, 11.76, 12.71, 12.13, _,
  _, _, _, _, _, _, _, 11.12, 7.62, 10.36, 11.08, 11.61, 11.82, 12.24, _,
  _, _, _, _, _, _, _, _, 9.33, 11.14, 11.62, 11.31, 12.1, 11.59, 11.67,
  _, _, _, _, _, _, _, _, 8.91, 11.79, 10.57, 12.02, 11.62, 11.51, _,
  _, _, _, _, _, _, _, _, _, 11.85, 9.66, 11.73, 11.21, _, _,
  _, _, _, _, _, _, _, _, _, 12, 10.52, 11.27, _, _, _,
  _, _, _, _, 10.46, 10.89, 11, _, _, 9.53, 9.05, 10.93, _, _, _,
  _, _, _, _, _, 10.43, _, 10.32, 9.25, 9.56, 9.45, _, _, _, _,
  _, _, _, _, _, _, _, 11.02, 9.7, 7.83, 9.97, _, _, _, _,
  _, _, _, _, _, _, _, 8.95, 9.23, 10.43, _, _, _, _, _,
  _, _, _, _, _, _, 8.86, 7.42, 8.62, 8.43, _, _, _, _, _,
  _, _, _, _, _, _, 10.45, 7.79, 6.97, 6.48, _, _, _, _, _,
  _, _, _, _, _, _, _, 6.88, 9.81, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 9.07, 7.94, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 13.98, _, 14.83, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 14.21, 14.65, 13.97, 15, 15.93, _, _, _,
  _, _, _, _, _, _, _, _, _, 15.4, 14.34, 14.68, 15.68, 15.1, _,
  _, _, _, _, _, _, _, 13.64, 10.02, 13.26, 14.01, 14.58, 14.81, 15.23, _,
  _, _, _, _, _, _, _, _, 11.88, 13.96, 14.45, 14.26, 15.05, 14.5, 14.63,
  _, _, _, _, _, _, _, _, 11.41, 14.49, 13.29, 14.95, 14.53, 14.34, _,
  _, _, _, _, _, _, _, _, _, 14.41, 12.19, 14.7, 14.2, _, _,
  _, _, _, _, _, _, _, _, _, 14.5, 13.23, 14.14, _, _, _,
  _, _, _, _, 13, 13.57, 13.58, _, _, 12.15, 11.89, 13.68, _, _, _,
  _, _, _, _, _, 13.01, _, 12.85, 11.87, 12.14, 12.2, _, _, _, _,
  _, _, _, _, _, _, _, 13.38, 12.23, 10.52, 12.64, _, _, _, _,
  _, _, _, _, _, _, _, 11.35, 11.67, 13.08, _, _, _, _, _,
  _, _, _, _, _, _, 10.91, 9.68, 11.29, 11.1, _, _, _, _, _,
  _, _, _, _, _, _, 12.53, 10.26, 9.7, 9.15, _, _, _, _, _,
  _, _, _, _, _, _, _, 9.17, 12.48, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 11.18, 10.36, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 15.97, _, 16.87, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 16.22, 16.66, 16.05, 17.13, 18.15, _, _, _,
  _, _, _, _, _, _, _, _, _, 17.36, 16.52, 16.98, 18.01, 17.62, _,
  _, _, _, _, _, _, _, 15.62, 12.1, 15.4, 16.29, 16.93, 17.26, 17.73, _,
  _, _, _, _, _, _, _, _, 13.87, 16.07, 16.61, 16.64, 17.48, 16.91, 17.19,
  _, _, _, _, _, _, _, _, 13.46, 16.52, 15.5, 17.23, 16.83, 16.79, _,
  _, _, _, _, _, _, _, _, _, 16.4, 14.25, 16.96, 16.64, _, _,
  _, _, _, _, _, _, _, _, _, 16.46, 15.31, 16.37, _, _, _,
  _, _, _, _, 14.74, 15.43, 15.48, _, _, 14.21, 14.2, 16.07, _, _, _,
  _, _, _, _, _, 14.85, _, 14.64, 13.76, 14.18, 14.45, _, _, _, _,
  _, _, _, _, _, _, _, 15.15, 14.19, 12.66, 14.98, _, _, _, _,
  _, _, _, _, _, _, _, 13.15, 13.56, 15.15, _, _, _, _, _,
  _, _, _, _, _, _, 12.74, 11.53, 13.29, 13.25, _, _, _, _, _,
  _, _, _, _, _, _, 14.33, 12.25, 11.97, 11.38, _, _, _, _, _,
  _, _, _, _, _, _, _, 11.16, 14.62, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 12.98, 12.48, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 16.26, _, 17.03, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 16.24, 16.5, 15.95, 16.93, 18.16, _, _, _,
  _, _, _, _, _, _, _, _, _, 17.16, 16.32, 16.74, 17.74, 17.49, _,
  _, _, _, _, _, _, _, 15.33, 11.99, 15.23, 15.96, 16.62, 17.07, 17.61, _,
  _, _, _, _, _, _, _, _, 13.6, 15.65, 16.35, 16.35, 17.36, 16.8, 17.11,
  _, _, _, _, _, _, _, _, 13.21, 16.29, 15.22, 17.03, 16.73, 16.84, _,
  _, _, _, _, _, _, _, _, _, 16.22, 14.03, 16.79, 16.5, _, _,
  _, _, _, _, _, _, _, _, _, 16.23, 14.9, 16.12, _, _, _,
  _, _, _, _, 14.45, 15.05, 15.3, _, _, 13.86, 13.86, 16.04, _, _, _,
  _, _, _, _, _, 14.54, _, 14.26, 13.44, 13.78, 14.17, _, _, _, _,
  _, _, _, _, _, _, _, 15.06, 13.83, 12.39, 14.82, _, _, _, _,
  _, _, _, _, _, _, _, 12.85, 13.31, 15.08, _, _, _, _, _,
  _, _, _, _, _, _, 12.61, 11.21, 12.89, 12.88, _, _, _, _, _,
  _, _, _, _, _, _, 14.13, 11.81, 11.53, 11.06, _, _, _, _, _,
  _, _, _, _, _, _, _, 10.97, 14.29, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 12.93, 12.24, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 14.77, _, 15.21, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 14.44, 14.32, 13.73, 14.43, 15.82, _, _, _,
  _, _, _, _, _, _, _, _, _, 14.75, 13.89, 14.16, 15.07, 14.86, _,
  _, _, _, _, _, _, _, 13.31, 10.01, 12.79, 13.44, 13.92, 14.41, 14.97, _,
  _, _, _, _, _, _, _, _, 11.47, 13.23, 13.82, 13.81, 14.79, 14.16, 14.56,
  _, _, _, _, _, _, _, _, 11.23, 13.96, 12.73, 14.45, 14.23, 14.51, _,
  _, _, _, _, _, _, _, _, _, 13.98, 11.72, 14.24, 14.04, _, _,
  _, _, _, _, _, _, _, _, _, 14.04, 12.54, 13.74, _, _, _,
  _, _, _, _, 12.37, 12.94, 13.37, _, _, 11.58, 11.46, 14.04, _, _, _,
  _, _, _, _, _, 12.53, _, 12.1, 11.25, 11.54, 11.9, _, _, _, _,
  _, _, _, _, _, _, _, 13.2, 11.48, 10.11, 12.62, _, _, _, _,
  _, _, _, _, _, _, _, 10.71, 11.03, 12.97, _, _, _, _, _,
  _, _, _, _, _, _, 10.74, 9.02, 10.39, 10.46, _, _, _, _, _,
  _, _, _, _, _, _, 12.19, 9.53, 9.12, 8.75, _, _, _, _, _,
  _, _, _, _, _, _, _, 8.86, 12.08, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 11.02, 10.07, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 12.27, _, 12.6, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 11.74, 11.19, 10.59, 11.2, 12.6, _, _, _,
  _, _, _, _, _, _, _, _, _, 11.4, 10.44, 10.77, 11.58, 11.39, _,
  _, _, _, _, _, _, _, 10.37, 7.02, 9.41, 10.01, 10.49, 10.84, 11.34, _,
  _, _, _, _, _, _, _, _, 8.55, 9.87, 10.32, 10.24, 11.18, 10.65, 10.95,
  _, _, _, _, _, _, _, _, 8.26, 10.66, 9.36, 10.89, 10.7, 11.13, _,
  _, _, _, _, _, _, _, _, _, 10.72, 8.51, 10.63, 10.49, _, _,
  _, _, _, _, _, _, _, _, _, 10.9, 9.23, 10.28, _, _, _,
  _, _, _, _, 9.43, 9.92, 10.48, _, _, 8.5, 8.19, 10.83, _, _, _,
  _, _, _, _, _, 9.59, _, 9.1, 8.17, 8.3, 8.8, _, _, _, _,
  _, _, _, _, _, _, _, 10.48, 8.25, 6.89, 9.47, _, _, _, _,
  _, _, _, _, _, _, _, 7.77, 7.82, 9.89, _, _, _, _, _,
  _, _, _, _, _, _, 8.06, 6.09, 7.1, 7.21, _, _, _, _, _,
  _, _, _, _, _, _, 9.5, 6.36, 5.92, 5.62, _, _, _, _, _,
  _, _, _, _, _, _, _, 5.96, 8.95, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 8.34, 7.16, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 9.61, _, 9.61, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 8.79, 7.93, 7.22, 7.6, 8.95, _, _, _,
  _, _, _, _, _, _, _, _, _, 7.89, 6.84, 7.07, 7.78, 7.62, _,
  _, _, _, _, _, _, _, 7.25, 4.07, 6.16, 6.38, 6.8, 6.98, 7.36, _,
  _, _, _, _, _, _, _, _, 5.5, 6.51, 6.76, 6.48, 7.2, 6.74, 6.9,
  _, _, _, _, _, _, _, _, 5.42, 7.28, 5.89, 7.2, 6.77, 7.32, _,
  _, _, _, _, _, _, _, _, _, 7.3, 5.12, 6.96, 6.66, _, _,
  _, _, _, _, _, _, _, _, _, 7.52, 5.92, 6.55, _, _, _,
  _, _, _, _, 6.43, 6.79, 7.55, _, _, 5.31, 4.97, 7.48, _, _, _,
  _, _, _, _, _, 6.63, _, 6.14, 5.13, 5.07, 5.57, _, _, _, _,
  _, _, _, _, _, _, _, 7.79, 5.05, 3.88, 6.16, _, _, _, _,
  _, _, _, _, _, _, _, 4.96, 4.78, 6.76, _, _, _, _, _,
  _, _, _, _, _, _, 5.46, 3.37, 4.02, 4.1, _, _, _, _, _,
  _, _, _, _, _, _, 6.87, 3.49, 2.93, 2.75, _, _, _, _, _,
  _, _, _, _, _, _, _, 3.13, 5.84, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 5.64, 4.15, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, 7.71, _, 7.42, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 6.64, 5.66, 4.9, 5.21, 6.35, _, _, _,
  _, _, _, _, _, _, _, _, _, 5.42, 4.41, 4.6, 5.36, 5.18, _,
  _, _, _, _, _, _, _, 5.08, 2.08, 3.91, 3.97, 4.32, 4.44, 4.82, _,
  _, _, _, _, _, _, _, _, 3.12, 4.07, 4.39, 3.94, 4.59, 4.15, 4.33,
  _, _, _, _, _, _, _, _, 3.25, 4.79, 3.47, 4.64, 4.21, 4.71, _,
  _, _, _, _, _, _, _, _, _, 4.77, 2.82, 4.43, 4.07, _, _,
  _, _, _, _, _, _, _, _, _, 4.98, 3.41, 3.98, _, _, _,
  _, _, _, _, 4.36, 4.78, 5.52, _, _, 2.85, 2.56, 5, _, _, _,
  _, _, _, _, _, 4.57, _, 3.94, 2.88, 2.62, 3.25, _, _, _, _,
  _, _, _, _, _, _, _, 5.59, 2.77, 1.58, 3.73, _, _, _, _,
  _, _, _, _, _, _, _, 2.87, 2.4, 4.28, _, _, _, _, _,
  _, _, _, _, _, _, 3.51, 1.22, 1.41, 1.77, _, _, _, _, _,
  _, _, _, _, _, _, 4.76, 1.3, 0.61, 0.53, _, _, _, _, _,
  _, _, _, _, _, _, _, 1, 3.41, _, _, _, _, _, _,
  _, _, _, _, _, _, _, 3.57, 1.92, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 transverse_mercator = _ ;

 latitude =
  47.844054553406, 47.8969525529387, 47.9443653984999, 47.9862574075524, 
    48.0225969129923, 48.0533563384176, 48.0785122641948, 48.0980454839399, 
    48.1119410510887, 48.1201883152932, 48.1227809484374, 48.1197169601269, 
    48.1109987025658, 48.0966328647939, 48.0766304563149,
  48.378619290464, 48.4325139474874, 48.4808218773753, 48.5235061454902, 
    48.5605339686372, 48.5918767947469, 48.6175103728438, 48.6374148128817, 
    48.651574635092, 48.6599788085598, 48.6626207788006, 48.659498484182, 
    48.6506143610939, 48.6359753378382, 48.6155928172742,
  48.9130218608792, 48.9679339810908, 49.0171557840908, 49.0606490234861, 
    49.0983797464768, 49.1303183782863, 49.156439796325, 49.1767233936352, 
    49.1911531312311, 49.1997175790201, 49.2024099450626, 49.1992280929964, 
    49.1901745475231, 49.1752564879247, 49.1544857296479,
  49.4472578366315, 49.5032090662785, 49.5533642947768, 49.5976839004742, 
    49.6361327039769, 49.6686800576857, 49.6952999244783, 49.7159709450422, 
    49.7306764934371, 49.739404720547, 49.7421485851522, 49.7389058724365, 
    49.7296791998144, 49.7144760100445, 49.6933085516707,
  49.9813225682174, 50.0383354373233, 50.0894444469083, 50.1346085324097, 
    50.1737912270996, 50.206960757122, 50.2340901250447, 50.255157181385, 
    50.2701446836498, 50.2790403425161, 50.2818368548624, 50.2785319234427, 
    50.2691282630822, 50.2536335933562, 50.2320606177962,
  50.5152111685507, 50.5733091369699, 50.6253931286521, 50.6714205639948, 
    50.7113536241457, 50.7451593519707, 50.7728097408599, 50.7942818107806, 
    50.809557671072, 50.8186245695759, 50.8214749277829, 50.8181063617693, 
    50.8085216887912, 50.7927289194921, 50.770741235776,
  51.0489184955607, 51.108126002083, 51.1612070673402, 51.208117519724, 
    51.2488181190882, 51.2832746641186, 51.3114580868158, 51.333344533439, 
    51.3489154313631, 51.3581575413985, 51.3610629952269, 51.3576293177042, 
    51.3478594338853, 51.3317616607229, 51.3093496834966,
  51.5824391333655, 51.6427816481124, 51.6968828169888, 51.7446967941835, 
    51.7861828443476, 51.8213054568834, 51.8500344465651, 51.8723450397762, 
    51.8882179457631, 51.8976394124096, 51.900601266152, 51.8971009357633, 
    51.8871414598433, 51.8707314779674, 51.8478852055503,
  52.1157673718818, 52.1772714522607, 52.2324167447687, 52.2811556415317, 
    52.3234458329554, 52.3592504295, 52.3885380689455, 52.411283008365, 
    52.4274652001427, 52.4370703514948, 52.4400899670742, 52.4365213743598, 
    52.4263677316542, 52.4096380186329, 52.386347009512,
  52.6488971847215, 52.7115905352255, 52.7678050163228, 52.8174911640789, 
    52.8606050100436, 52.8971082111323, 52.9269681640948, 52.9501581037095, 
    52.9666571839719, 52.9764505416834, 52.979529341976, 52.9758908054466, 
    52.965538216704, 52.9484809142686, 52.9247342618969,
  53.1818222052031, 53.2457337413763, 53.3030435798176, 53.3537002998775, 
    53.3976581835935, 53.4348773543624, 53.465323899227, 53.4889699738255, 
    53.5057938891998, 53.5157801798047, 53.5189196522095, 53.5152094141286, 
    53.5046528835675, 53.4872597780149, 53.4630460837632,
  53.7145357002922, 53.7796956172061, 53.8381281485985, 53.8897798092197, 
    53.9346030343673, 53.9725563281028, 54.0036043940333, 54.0277182476074, 
    54.0448753090365, 54.0550594761175, 54.0582611763918, 54.054477398243, 
    54.0437117006932, 54.0259742018267, 54.0012815459257,
  54.2470305422583, 54.3134703878825, 54.373054182306, 54.4257262599315, 
    54.4714371049381, 54.5101435098718, 54.5418087156705, 54.5664025319582, 
    54.5839014366276, 54.5942886539082, 54.5975542102961, 54.5936949679049, 
    54.5827146349733, 54.564623753448, 54.5394396637395,
  54.7792991778142, 54.8470519317006, 54.9078168662906, 54.9615360113346, 
    55.0081577877224, 55.0476371773658, 55.0799358732922, 55.1050224086606, 
    55.1228722636109, 55.1334679490571, 55.1367990667356, 55.1328623450157, 
    55.1216616501845, 55.1032079731123, 55.0775193914075,
  55.3113335944753, 55.3804337522171, 55.4424110891485, 55.4972051967358, 
    55.5447623119092, 55.5850354992511, 55.6179848120742, 55.6435774309587, 
    55.6617877785416, 55.6725976095683, 55.6759960754424, 55.6719797627292, 
    55.6605527052888, 55.641726369938, 55.615519615762,
  55.843125283842, 55.9136089478164, 55.9768314181721, 56.0327297042825, 
    56.081247729164, 56.1223365250921, 56.1559544066787, 56.1820671198206, 
    56.2006479651745, 56.21167789506, 56.2151455829404, 56.2110474648736, 
    56.1993877525764, 56.1801784179872, 56.1534391494615,
  56.3746652014777, 56.4465701784313, 56.51107207249, 56.5681051560061, 
    56.6176108979737, 56.6595381743173, 56.693843454095, 56.7204909598463, 
    56.7394528005849, 56.7507090762136, 56.754247952412, 56.750065705323, 
    56.7381667356373, 56.71856355195, 56.6912767235385,
  56.9059437230068, 56.9793096291045, 57.0451268936382, 57.103326884848, 
    57.1538484664777, 57.196638224117, 57.2316506657855, 57.2588483947802, 
    57.2782022531129, 57.2896914341739, 57.29330356356, 57.2890347473156, 
    57.2768895871385, 57.2568811624115, 57.2290309792247,
  57.4369505960174, 57.5118189700359, 57.578989313273, 57.6383899094422, 
    57.6899568536137, 57.7336342961484, 57.7693746590588, 57.7971388225841, 
    57.816896280109, 57.8286252598986, 57.832312812463, 57.8279548627103, 
    57.8155562263881, 57.7951305906551, 57.7667004589706,
  57.9676748872937, 58.0440893127173, 58.1126523176974, 58.1732889063911, 
    58.2259322283806, 58.2705238419087, 58.3070139475765, 58.3353615900183, 
    58.3555348254607, 58.3675108534508, 58.3712761114255, 58.3668263311779, 
    58.3541665566602, 58.3333111229464, 58.3042835965647,
  58.498104924846, 58.5761111617035, 58.6461084088293, 58.7080181797435, 
    58.7617704869969, 58.8073041266193, 58.8445669308941, 58.8735159866727, 
    58.8941178168711, 58.9063485232267, 58.9101938888227, 58.9056494393177, 
    58.8927204622524, 58.8714219842362, 58.8417787062455,
  59.0282282341341, 59.1078743615042, 59.1793495611899, 59.2425716273373, 
    59.2974672277007, 59.3439722114381, 59.3820318829152, 59.411601238381, 
    59.4326451628626, 59.4451385851145, 59.4490665889397, 59.4444244796915, 
    59.4312178052443, 59.4094623312131, 59.3791839706838,
  59.5580314677991, 59.6393680380188, 59.7123671744334, 59.7769427036279, 
    59.8330177229016, 59.8805249337978, 59.919406939127, 59.9496164999416, 
    59.9711167494711, 59.9838813615732, 59.9878946718049, 59.983151749767, 
    59.9696584219201, 59.9474312446241, 59.9164974276951,
  60.0875003281259, 60.1705805338489, 60.2451520208694, 60.311124378567, 
    60.3684168883567, 60.4169588856313, 60.4566900824628, 60.487560847059, 
    60.5095324365905, 60.5225771806242, 60.5266786130184, 60.5218315507563, 
    60.5080421188128, 60.485327720771, 60.4537169555242,
  60.6166194813516, 60.7014993367357, 60.7776941873556, 60.8451090920328, 
    60.9036592489909, 60.9532703892175, 60.9938791276155, 61.0254332674031, 
    61.0478920539255, 61.0612263747446, 61.0654189035752, 61.0604641863409, 
    61.0463686683224, 61.023150662078, 60.990840256516 ;

 longitude =
  -9.98920028497714, -9.19383379941614, -8.39629883287295, -7.59682698288458, 
    -6.7956534930323, -5.99301683616649, -5.18915828099242, 
    -4.38432144440827, -3.5787518319865, -2.77269636898997, 
    -1.96640292431389, -1.16011982974503, -0.354095396929169, 
    0.451422565561637, 1.25618723267107,
  -10.0730473274966, -9.26952262947054, -8.46374772716654, -7.65596265450841, 
    -6.84641132860804, -6.03534110711392, -5.22300232734314, 
    -4.40964782981475, -3.59553246880245, -2.78091261252458, 
    -1.96604563558933, -1.15118940631312, -0.336601771530144, 
    0.477459958489061, 1.29073952239195,
  -10.1593810431334, -9.34746236100672, -8.53320743066179, -7.71686514993805, 
    -6.89868855574897, -6.07893435363003, -5.25786242731941, 
    -4.43573533124081, -3.61281776875803, -2.78937605907095, 
    -1.96567759562231, -1.14199029888498, -0.318582066399204, 
    0.50427977707058, 1.32632902638977,
  -10.2482961032679, -9.42773908227278, -8.60475516492533, -7.77960256701633, 
    -6.95254391977765, -6.12384576954099, -5.29377805548334, 
    -4.46261356860862, -3.63062739511449, -2.7980963472936, 
    -1.96529838511857, -1.13251203165965, -0.30001578548457, 
    0.531912466810522, 1.36299603478965,
  -10.3398922183497, -9.51044348905737, -8.67847230493588, -7.84424668223468, 
    -7.00803935141737, -6.17012722466197, -5.33079083928247, 
    -4.49031378053214, -3.64898208724899, -2.80708364380385, 
    -1.9649075618113, -1.12274355506411, -0.280881311151358, 
    0.560390136779237, 1.40078303465438,
  -10.4342744706801, -9.59567119112506, -8.75444465705699, -7.91087319829539, 
    -7.06524018218587, -6.21783344647522, -5.36894470569428, 
    -4.51886893485574, -3.66790373427435, -2.81634867931662, 
    -1.96450465888738, -1.11267320646047, -0.261155827460731, 
    0.589746673195278, 1.43973485959274,
  -10.5315536738368, -9.68352304339319, -8.83276275962293, -7.97956201194649, 
    -7.12421537752807, -6.267022216842, -5.40828604005279, -4.54831384840343, 
    -3.68741545480617, -2.82590278783039, -1.9640891832819, 
    -1.10228866756811, -0.240815237043595, 0.620017862469661, 1.47989885179272,
  -10.6318467612406, -9.77410550419627, -8.91352220830109, -8.05039750404384, 
    -7.18503778940964, -6.31775458521625, -5.44886385825236, 
    -4.57868531684511, -3.70754168348402, -2.83575794912879, 
    -1.96366061382805, -1.09157691827639, -0.21983407093693, 
    0.651241524643249, 1.52132503769771,
  -10.7352772066352, -9.86753102323976, -8.99682400863316, -8.12346885401316, 
    -7.2477844302867, -6.37009509999337, -5.49072999365883, 
    -4.61002225568976, -3.72830826492246, -2.84592683493686, 
    -1.96321839924786, -1.0805241864859, -0.198185390678629, 
    0.683457658254388, 1.56406631868217,
  -10.8419754795513, -9.96391846213299, -9.0827749584256, -8.19887038112937, 
    -7.31253677058499, -6.42411205981478, -5.53393930021181, 
    -4.64236585353224, -3.74974255584634, -2.85642285910366, 
    -1.96276195596758, -1.06911589357479, -0.175840681874954, 
    0.716708597793942, 1.60817867823921,
  -10.9520795391697, -10.063393550715, -9.17148806296315, -8.27670191530788, 
    -7.37938106206783, -6.47987778686049, -5.57854987337538, 
    -4.67575973881273, -3.77187353625348, -2.86726023222659, 
    -1.96229066573964, -1.0573365950385, -0.152769738362318, 
    0.751039185040595, 1.65372140736972,
  -11.0657353703763, -10.1660893827517, -9.26308298636029, -8.35706920041487, 
    -7.44840868975096, -6.53746892440155, -5.6246232907905, 
    -4.71025016149765, -3.79473193054869, -2.87845402118278, 
    -1.96180387305082, -1.04516991579751, -0.128940535980074, 
    0.786496955723276, 1.7007573500622,
  -11.1830975662371, -10.2721469549954, -9.3576865427521, -8.44008433345767, 
    -7.51971655533774, -6.59696676115596, -5.67222487470614, 
    -4.74588619126134, -3.8183503397075, -2.89002021408905, 
    -1.96130088229406, -1.0325984796063, -0.104319094851846, 
    0.82313234313237, 1.74935317098051,
  -11.3043299616042, -10.381715754062, -9.45543323146308, -8.52586624341769, 
    -7.59340749550684, -6.65845758530051, -5.72142397851931, 
    -4.78271993394163, -3.84276338565827, -2.90197579127684, 
    -1.96078095467818, -1.01960383192669, -0.0788693289371003, 
    0.860998900500445, 1.7995796477347,
  -11.4296063231135, -10.4949543961106, -9.55646582078833, -8.61454121394411, 
    -7.66959073879178, -6.72203307134266, -5.77229430004354, 
    -4.82080676826331, -3.86800786922023, -2.91433880294146, 
    -1.96024330484687, -1.00616635554885, -0.052552881459902, 
    0.900153544200024, 1.85151199040478,
  -11.5591111014597, -10.6120313249043, -9.66093598558494, -8.7062434546453, 
    -7.74838240525585, -6.78779070345745, -5.82491422445522, 
    -4.86020560507619, -3.89412294310471, -2.9271284542093, 
    -1.95968709717459, -0.992265178152314, -0.0253289446447839, 
    0.94065682006507, 1.90523019132359,
  -11.6930402525323, -10.7331255745149, -9.76900500451231, -8.80111572630578, 
    -7.82990605369611, -6.85583423935267, -5.87936720024468, 
    -4.90097917164317, -3.92115030168147, -2.94036519846278, 
    -1.9591114417026, -0.977878070894472, 0.00284593801297501, 
    0.982573195439496, 1.960819408509,
  -11.8316021348019, -10.8584276037011, -9.88084452349077, -8.8993100260318, 
    -7.91429328171586, -6.92627421925024, -5.93574215193132, 
    -4.94319432384538, -3.9491343894355, -2.9540708398732, -1.95851538967384, 
    -0.962981336994358, 0.0320180889478738, 1.02597137989613, 2.01837038657676,
  -11.9750184912516, -10.9881402098746, -9.99663739278248, -9.0009883391005, 
    -8.00168438469909, -6.99922852517364, -5.99413393379908, 
    -4.98692238955231, -3.97812263029623, -2.96826864621866, 
    -1.95789792861975, -0.947549689141366, 0.0622369354681829, 
    1.07092467796048, 2.07797991947095,
  -12.1235255251842, -11.1224795315696, -10.1165785860531, -9.10632346517315, 
    -8.0922290805179, -7.07482299642293, -6.05464382948011, 
    -5.03223954684354, -4.00816568031739, -2.98298347321084, 
    -1.9572579769454, -0.9315561143995, 0.0935552730242402, 1.11751137762407, 
    2.13975135993129,
  -12.2773750804151, -11.2616761494831, -10.2408762108673, -9.21549992754912, 
    -8.18608730772077, -7.15319210791668, -6.11738010287401, 
    -5.07922724127552, -4.03931770652723, -2.99824190172356, 
    -1.95659437795255, -0.914971725093862, 0.126029555737895, 
    1.16581517895175, 2.20379518128831,
  -12.4368359377125, -11.4059762974686, -10.3697526213277, -9.32871497530801, 
    -8.28343010600673, -7.2344797190002, -6.18245860665242, 
    -5.12797264697275, -4.07163669516534, -3.01407238951204, 
    -1.95590589323104, -0.897765593953164, 0.15972021754213, 
    1.21592566768898, 2.27022959795357,
  -12.6021952408859, -11.5556431963767, -10.5034456450135, -9.4461796895363, 
    -8.38444058901275, -7.31883990138514, -6.25000345548213, 
    -5.17856917700279, -4.10518479298119, -3.03050543923978, 
    -1.95519119533947, -0.879904571534727, 0.194692027758326, 
    1.26793883947262, 2.33918125187156,
  -12.7737600676953, -11.7109585253746, -10.642209938044, -9.56812020639526, 
    -8.48931502085637, -7.4064378561215, -6.32014777212634, 
    -5.23111704928498, -4.14002868580464, -3.0475737848944, 
    -1.95444885968423, -0.861353083670598, 0.231014485495231, 
    1.3219576810598, 2.41078597324487,
  -12.9518591627846, -11.8722240473793, -10.7863184840172, -9.69477907159376, 
    -8.59826400951848, -7.49745093094017, -6.39303451577815, 
    -5.28572391520457, -4.17624001922245, -3.06531259898384, 
    -1.95367735549274, -0.842072906337468, 0.268762257903138, 
    1.3780928159349, 2.48518962506041 ;

 projection_x_coordinate = -197500, -137500, -77500, -17500, 42500, 102500, 
    162500, 222500, 282500, 342500, 402500, 462500, 522500, 582500, 642500 ;

 projection_x_coordinate_bnds =
  -200000, -195000,
  -140000, -135000,
  -80000, -75000,
  -20000, -15000,
  40000, 45000,
  100000, 105000,
  160000, 165000,
  220000, 225000,
  280000, 285000,
  340000, 345000,
  400000, 405000,
  460000, 465000,
  520000, 525000,
  580000, 585000,
  640000, 645000 ;

 projection_y_coordinate = -197500, -137500, -77500, -17500, 42500, 102500, 
    162500, 222500, 282500, 342500, 402500, 462500, 522500, 582500, 642500, 
    702500, 762500, 822500, 882500, 942500, 1002500, 1062500, 1122500, 
    1182500, 1242500 ;

 projection_y_coordinate_bnds =
  -200000, -195000,
  -140000, -135000,
  -80000, -75000,
  -20000, -15000,
  40000, 45000,
  100000, 105000,
  160000, 165000,
  220000, 225000,
  280000, 285000,
  340000, 345000,
  400000, 405000,
  460000, 465000,
  520000, 525000,
  580000, 585000,
  640000, 645000,
  700000, 705000,
  760000, 765000,
  820000, 825000,
  880000, 885000,
  940000, 945000,
  1000000, 1005000,
  1060000, 1065000,
  1120000, 1125000,
  1180000, 1185000,
  1240000, 1245000 ;

 time = 1586976, 1587720, 1588392, 1589136, 1589856, 1590600, 1591320, 
    1592064, 1592808, 1593528, 1594272, 1594992 ;

 season_year = 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;
}
